magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 612 108 648
rect 0 576 144 612
rect 0 540 180 576
rect 36 504 216 540
rect 72 468 252 504
rect 108 432 288 468
rect 144 324 324 432
rect 108 288 288 324
rect 72 252 252 288
rect 36 216 216 252
rect 0 180 180 216
rect 0 144 144 180
rect 0 108 108 144
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
