VERSION 5.8 ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS
        
LAYER M2
    TYPE ROUTING ;
    WIDTH 0.2 ;
END M2

END LIBRARY
