* Extracted by KLayout

* cell TOP
* pin A
* pin C
* pin SUBSTRATE
.SUBCKT TOP 2 3 4
* net 2 A
* net 3 C
* net 4 SUBSTRATE
* cell instance $1 r0 *1 0,0
X$1 2 3 1 6 4 DINV
* cell instance $2 r0 *1 3.6,0
X$2 5 6 1 4 INVX1
.ENDS TOP

* cell DINV
* pin A<1>
* pin A<2>
* pin B<2>
* pin VDD
* pin VSS
.SUBCKT DINV 1 2 3 5 6
* net 1 A<1>
* net 2 A<2>
* net 3 B<2>
* net 4 B<1>
* net 5 VDD
* net 6 VSS
* cell instance $1 r0 *1 0,0
X$1 4 5 1 6 INVX1
* cell instance $2 r0 *1 1.8,0
X$2 3 5 2 6 INVX1
.ENDS DINV

* cell INVX1
* pin OUT
* pin VDD
* pin IN
* pin VSS
.SUBCKT INVX1 1 2 3 4
* net 1 OUT
* net 2 VDD
* net 3 IN
* net 4 VSS
* device instance $1 r0 *1 0.85,2.135 NMOS
M$1 4 3 1 4 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $2 r0 *1 0.85,5.8 PMOS
M$2 2 3 1 2 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
.ENDS INVX1
