* written by unit test

* cell SUBCKT
* pin 
* pin A
* pin V42
* pin Z
* pin gnd
* pin gnd
.SUBCKT SUBCKT \$1 A[5]<1> V42\x28\x25\x29 Z gnd gnd$1
XD_$1 V42\x28\x25\x29 \$3 Z \$1 HVPMOS PARAMS: L=0.2 W=1 AS=0.18 AD=0.18
+ PS=2.16 PD=2.16
* device instance $2 r0 *1 0,0 HVPMOS
XD_$2 V42\x28\x25\x29 A[5]<1> \$3 \$1 HVPMOS PARAMS: L=0.2 W=1 AS=0.18 AD=0.18
+ PS=2.16 PD=2.16
XD_$3 gnd \$3 gnd gnd$1 HVNMOS PARAMS: L=1.13 W=2.12 PS=6 PD=6 AS=0 AD=0
XD_$4 gnd \$3 Z gnd$1 HVNMOS PARAMS: L=0.4 W=0.4 PS=1.16 PD=1.16 AS=0.19 AD=0.19
XD_$5 gnd A[5]<1> \$3 gnd$1 HVNMOS PARAMS: L=0.4 W=0.4 PS=1.76 PD=1.76 AS=0.19 AD=0.19
.ENDS SUBCKT
.SUBCKT SUBCKT \$1 A[5]<1> V42\x28\x25\x29 Z gnd gnd$1
XD_$13 gnd \$3 gnd gnd$1 HVNMOS PARAMS: L=1.13 W=2.12 PS=6 PD=6 AS=0 AD=0
.ENDS SUBCKT
