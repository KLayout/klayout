magic
tech scmos
timestamp 1534344057
<< silk >>
rect 2 17 12 18
rect 1 16 12 17
rect 0 14 12 16
rect 0 10 4 14
rect 0 6 10 10
rect 0 0 4 6
<< end >>
