magic
tech scmos
timestamp 1543784536
use Library/magic/L500_CHAR_u  L500_CHAR_u_0
timestamp 1534323899
transform 1 0 20 0 1 272
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_4
timestamp 1534321786
transform 1 0 36 0 1 272
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_2
timestamp 1534323853
transform 1 0 52 0 1 280
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_3
timestamp 1534323853
transform 1 0 68 0 1 280
box 0 0 12 18
use Library/magic/L500_CHAR_g  L500_CHAR_g_0
timestamp 1534322005
transform 1 0 4 0 1 268
box 0 0 12 18
use Library/magic/T7_INV  T7_INV_0
timestamp 1533657739
transform 1 0 0 0 1 188
box 0 0 16 56
use Library/magic/T10_NAND2  T10_NAND2_0
timestamp 1533654735
transform 1 0 26 0 1 188
box 0 0 24 80
use Library/magic/T11_NOR2  T11_NOR2_0
timestamp 1533654819
transform 1 0 60 0 1 188
box 0 0 24 88
use Library/magic/L500_CHAR_a  L500_CHAR_a_1
timestamp 1534325357
transform 1 0 130 0 1 274
box 0 0 12 18
use Library/magic/L500_CHAR_t  L500_CHAR_t_0
timestamp 1534318840
transform 1 0 146 0 1 274
box 0 0 12 18
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_3
timestamp 1534325697
transform 1 0 166 0 1 282
box 0 0 4 4
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_4
timestamp 1534325697
transform 1 0 174 0 1 282
box 0 0 4 4
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_5
timestamp 1534325697
transform 1 0 182 0 1 282
box 0 0 4 4
use Library/magic/L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 94 0 1 268
box 0 0 16 18
use Library/magic/L500_CHAR_h  L500_CHAR_h_0
timestamp 1534224731
transform 1 0 114 0 1 268
box 0 0 12 18
use Library/magic/T7_NAND2  T7_NAND2_0
timestamp 1533654698
transform 1 0 94 0 1 188
box 0 0 24 56
use Library/magic/T10_NAND3  T10_NAND3
timestamp 1533654785
transform 1 0 128 0 1 188
box 0 0 32 80
use Library/magic/T11_NOR3  T11_NOR3_0
timestamp 1533654861
transform 1 0 170 0 1 188
box 0 0 32 88
use Library/magic/L500_CHAR_l  L500_CHAR_l_1
timestamp 1534225390
transform 1 0 8 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 24 0 1 164
box 0 0 8 18
use Library/magic/L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 36 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_r  L500_CHAR_r_1
timestamp 1534323573
transform 1 0 52 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_3
timestamp 1534321786
transform 1 0 68 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_1
timestamp 1534323853
transform 1 0 88 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_1
timestamp 1534226087
transform 1 0 104 0 1 164
box 0 0 8 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_2
timestamp 1534225390
transform 1 0 116 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_2
timestamp 1534226087
transform 1 0 132 0 1 164
box 0 0 8 18
use Library/magic/L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 144 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_o  L500_CHAR_o_0
timestamp 1534323159
transform 1 0 160 0 1 164
box 0 0 12 18
use Library/magic/L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 176 0 1 164
box 0 0 12 18
use Library/magic/L500_SIGNATURE_pearlriver  L500_SIGNATURE_pearlriver_0
timestamp 1543784536
transform 1 0 0 0 1 142
box 0 0 202 18
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_0
timestamp 1534325697
transform 1 0 16 0 1 120
box 0 0 4 4
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_1
timestamp 1534325697
transform 1 0 24 0 1 120
box 0 0 4 4
use Library/magic/L500_CHAR_dot  L500_CHAR_dot_2
timestamp 1534325697
transform 1 0 32 0 1 120
box 0 0 4 4
use Library/magic/L500_CHAR_r  L500_CHAR_r_0
timestamp 1534323573
transform 1 0 44 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 60 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 76 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_1
timestamp 1534321786
transform 1 0 92 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 108 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_s  L500_CHAR_s_0
timestamp 1534323853
transform 1 0 124 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_2
timestamp 1534321786
transform 1 0 140 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 156 0 1 120
box 0 0 12 18
use Library/magic/L500_CHAR_mark  L500_CHAR_mark_0
timestamp 1534327094
transform 1 0 172 0 1 120
box 0 0 4 18
use Library/magic/L500_SIGNATURE_kallisti  L500_SIGNATURE_kallisti_0
timestamp 1533657739
transform 1 0 40 0 1 -4
box 4 4 116 118
<< end >>
