* Tests the ability to translate subcircuits into plain devices

.SUBCKT HVNMOS S G D B PARAMS: L=0 W=0 AS=0 AD=0 PS=0 PD=0
MINT S G D B MODEL L=L W=W AS=AS AD=AD PS=PS PD=PD
* parasitic stuff
C1 S G 1.5F*L+5.5*L*W
C2 D G 1.2F*L+5.5*L*W
C3 S B 2.1F*AS+0.2*PS
C4 D B 2.1F*AD+0.2*PD
.ENDS HVNMOS

.SUBCKT HVPMOS S G D B PARAMS: L=0 W=0 AS=0 AD=0 PS=0 PD=0
MINT S G D B MODEL L=L W=W AS=AS AD=AD
* parasitic stuff
C1 S G 0.8F*L+4.2*L*W
C2 D G 0.8F*L+4.2*L*W
C3 S B 2.5F*AS+0.3*PS
C4 D B 2.5F*AD+0.3*PD
.ENDS HVPMOS

.SUBCKT SUBCKT \$1 A VDD Z gnd gnd$1
X$1 VDD \$3 Z \$1 HVPMOS PARAMS: L=0.2 W=1 AS=0.18 AD=0.18 PS=2.16 PD=2.16
X$2 VDD A \$3 \$1 HVPMOS PARAMS: L=0.2 W=1 AS=0.18 AD=0.18 PS=2.16 PD=2.16
X$3 gnd \$3 gnd gnd$1 HVNMOS PARAMS: L=1.13 W=2.12 PS=6 PD=6 AS=0 AD=0
X$4 gnd \$3 Z gnd$1 HVNMOS PARAMS: L=0.4 W=0.4 PS=1.16 PD=1.16 AS=0.19 AD=0.19
X$5 gnd A \$3 gnd$1 HVNMOS PARAMS: L=0.4 W=0.4 PS=1.76 PD=1.76 AS=0.19 AD=0.19
.ENDS SUBCKT

XSUBCKT IN OUT VDD Z VSS VSS SUBCKT

