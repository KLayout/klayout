* Extracted by KLayout

.SUBCKT TOP A Q VDD SUBSTRATE|VSS
X$1 SUBSTRATE|VSS VDD \$1 Q INV
X$2 SUBSTRATE|VSS VDD A \$1 INV
.ENDS TOP

.SUBCKT INV SUBSTRATE \$2 \$4 \$5
M$1 \$2 \$4 \$5 \$2 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
M$2 SUBSTRATE \$4 \$5 SUBSTRATE NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P
+ PS=3.45U PD=3.45U
.ENDS INV
