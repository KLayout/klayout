magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 108 540 216 756
rect 324 540 432 756
rect 0 432 540 540
rect 108 324 216 432
rect 324 324 432 432
rect 0 216 540 324
rect 108 0 216 216
rect 324 0 432 216
<< properties >>
string FIXED_BBOX 0 -216 648 756
<< end >>
