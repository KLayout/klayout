magic
timestamp 1575832387
<< checkpaint >>
rect -1 0 25 80
<< l5d0 >>
rect 14 29 17 48
rect 7 29 10 48
<< l1001d0 >>
rect 0 20 24 24
rect 0 29 24 33
rect 0 38 24 42
rect 0 47 24 51
rect 0 56 24 60
<< l8d0 >>
rect 18 63 20 64
rect 18 52 20 53
rect 18 57 20 59
rect 4 63 6 64
rect 4 57 6 59
rect 11 52 13 53
rect 4 52 6 53
rect 11 63 13 64
rect 11 57 13 59
rect 18 18 20 20
rect 4 18 6 20
rect 18 23 20 25
rect 4 23 6 25
<< l9d0 >>
rect 18 17 21 28
rect 18 28 22 31
rect 19 31 22 45
rect 4 45 22 48
rect 4 48 7 51
rect 0 4 24 12
rect 0 68 24 76
rect 18 51 21 65
rect 4 51 7 65
rect 11 51 14 68
rect 18 48 21 51
rect 4 12 7 26
<< l13d0 >>
rect 0 0 24 80
<< l1d0 >>
rect -1 45 25 80
<< l14d0 >>
rect 9 49 16 67
rect 9 13 16 28
<< labels >>
rlabel l9d0 12.5 72 12.5 72 0 VDD
rlabel l9d0 12.5 8 12.5 8 0 VSS
rlabel l9d0 21 40 21 40 0 OUT
rlabel l9d0 8 31 8 31 0 A
rlabel l9d0 15 40 15 40 0 B
use POLYM1 POLYM1_1
timestamp 1575832387
transform 1 0 8 0 1 31
box -5 -5 5 5
use POLYM1 POLYM1_2
timestamp 1575832387
transform 1 0 15 0 1 40
box -5 -5 5 5
use NMOS2 NMOS2_1
timestamp 1575832387
transform 1 0 3 0 1 17
box -1 -3 12 12
use PMOS3 PMOS3_1
timestamp 1575832387
transform 1 0 3 0 1 51
box -1 -3 12 18
use PMOS3 PMOS3_2
timestamp 1575832387
transform 1 0 10 0 1 51
box -1 -3 12 18
use NMOS2 NMOS2_2
timestamp 1575832387
transform 1 0 10 0 1 17
box -1 -3 12 12
<< end >>
