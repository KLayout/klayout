magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 396 108 756
rect 216 396 324 756
rect 0 324 324 396
rect 36 216 288 324
rect 72 108 252 216
rect 108 0 216 108
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
