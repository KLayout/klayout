magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 0 432 108
<< properties >>
string FIXED_BBOX 0 -216 540 756
<< end >>
