magic
tech scmos
timestamp 1533657739
<< silk >>
rect 182 234 183 235
rect 183 234 184 235
rect 181 233 182 234
rect 182 233 183 234
rect 183 233 184 234
rect 184 233 185 234
rect 185 233 186 234
rect 180 232 181 233
rect 181 232 182 233
rect 182 232 183 233
rect 183 232 184 233
rect 184 232 185 233
rect 185 232 186 233
rect 179 231 180 232
rect 180 231 181 232
rect 181 231 182 232
rect 182 231 183 232
rect 183 231 184 232
rect 184 231 185 232
rect 185 231 186 232
rect 177 230 178 231
rect 178 230 179 231
rect 179 230 180 231
rect 180 230 181 231
rect 181 230 182 231
rect 182 230 183 231
rect 183 230 184 231
rect 184 230 185 231
rect 185 230 186 231
rect 186 230 187 231
rect 176 229 177 230
rect 177 229 178 230
rect 178 229 179 230
rect 179 229 180 230
rect 180 229 181 230
rect 181 229 182 230
rect 182 229 183 230
rect 183 229 184 230
rect 184 229 185 230
rect 185 229 186 230
rect 186 229 187 230
rect 187 229 188 230
rect 176 228 177 229
rect 177 228 178 229
rect 178 228 179 229
rect 179 228 180 229
rect 180 228 181 229
rect 181 228 182 229
rect 182 228 183 229
rect 183 228 184 229
rect 184 228 185 229
rect 185 228 186 229
rect 186 228 187 229
rect 187 228 188 229
rect 176 227 177 228
rect 177 227 178 228
rect 178 227 179 228
rect 179 227 180 228
rect 180 227 181 228
rect 181 227 182 228
rect 182 227 183 228
rect 183 227 184 228
rect 184 227 185 228
rect 185 227 186 228
rect 186 227 187 228
rect 187 227 188 228
rect 175 226 176 227
rect 176 226 177 227
rect 177 226 178 227
rect 178 226 179 227
rect 179 226 180 227
rect 180 226 181 227
rect 181 226 182 227
rect 182 226 183 227
rect 183 226 184 227
rect 184 226 185 227
rect 185 226 186 227
rect 186 226 187 227
rect 187 226 188 227
rect 188 226 189 227
rect 174 225 175 226
rect 175 225 176 226
rect 176 225 177 226
rect 177 225 178 226
rect 178 225 179 226
rect 179 225 180 226
rect 180 225 181 226
rect 181 225 182 226
rect 182 225 183 226
rect 183 225 184 226
rect 184 225 185 226
rect 185 225 186 226
rect 186 225 187 226
rect 187 225 188 226
rect 188 225 189 226
rect 173 224 174 225
rect 174 224 175 225
rect 175 224 176 225
rect 176 224 177 225
rect 177 224 178 225
rect 178 224 179 225
rect 179 224 180 225
rect 180 224 181 225
rect 181 224 182 225
rect 182 224 183 225
rect 183 224 184 225
rect 184 224 185 225
rect 185 224 186 225
rect 186 224 187 225
rect 187 224 188 225
rect 188 224 189 225
rect 172 223 173 224
rect 173 223 174 224
rect 174 223 175 224
rect 175 223 176 224
rect 176 223 177 224
rect 177 223 178 224
rect 178 223 179 224
rect 179 223 180 224
rect 180 223 181 224
rect 181 223 182 224
rect 182 223 183 224
rect 183 223 184 224
rect 184 223 185 224
rect 185 223 186 224
rect 186 223 187 224
rect 187 223 188 224
rect 188 223 189 224
rect 189 223 190 224
rect 172 222 173 223
rect 173 222 174 223
rect 174 222 175 223
rect 175 222 176 223
rect 176 222 177 223
rect 177 222 178 223
rect 178 222 179 223
rect 179 222 180 223
rect 180 222 181 223
rect 181 222 182 223
rect 182 222 183 223
rect 183 222 184 223
rect 184 222 185 223
rect 185 222 186 223
rect 186 222 187 223
rect 187 222 188 223
rect 188 222 189 223
rect 189 222 190 223
rect 171 221 172 222
rect 172 221 173 222
rect 173 221 174 222
rect 174 221 175 222
rect 175 221 176 222
rect 176 221 177 222
rect 177 221 178 222
rect 178 221 179 222
rect 179 221 180 222
rect 180 221 181 222
rect 181 221 182 222
rect 182 221 183 222
rect 183 221 184 222
rect 184 221 185 222
rect 185 221 186 222
rect 186 221 187 222
rect 187 221 188 222
rect 188 221 189 222
rect 189 221 190 222
rect 170 220 171 221
rect 171 220 172 221
rect 172 220 173 221
rect 173 220 174 221
rect 174 220 175 221
rect 175 220 176 221
rect 176 220 177 221
rect 177 220 178 221
rect 178 220 179 221
rect 179 220 180 221
rect 180 220 181 221
rect 181 220 182 221
rect 182 220 183 221
rect 183 220 184 221
rect 184 220 185 221
rect 185 220 186 221
rect 186 220 187 221
rect 187 220 188 221
rect 188 220 189 221
rect 189 220 190 221
rect 169 219 170 220
rect 170 219 171 220
rect 171 219 172 220
rect 172 219 173 220
rect 173 219 174 220
rect 174 219 175 220
rect 175 219 176 220
rect 176 219 177 220
rect 177 219 178 220
rect 178 219 179 220
rect 179 219 180 220
rect 180 219 181 220
rect 181 219 182 220
rect 182 219 183 220
rect 183 219 184 220
rect 184 219 185 220
rect 185 219 186 220
rect 186 219 187 220
rect 187 219 188 220
rect 188 219 189 220
rect 189 219 190 220
rect 112 218 113 219
rect 113 218 114 219
rect 114 218 115 219
rect 115 218 116 219
rect 116 218 117 219
rect 117 218 118 219
rect 118 218 119 219
rect 119 218 120 219
rect 120 218 121 219
rect 121 218 122 219
rect 122 218 123 219
rect 168 218 169 219
rect 169 218 170 219
rect 170 218 171 219
rect 171 218 172 219
rect 172 218 173 219
rect 173 218 174 219
rect 174 218 175 219
rect 175 218 176 219
rect 176 218 177 219
rect 177 218 178 219
rect 178 218 179 219
rect 179 218 180 219
rect 180 218 181 219
rect 181 218 182 219
rect 182 218 183 219
rect 183 218 184 219
rect 184 218 185 219
rect 185 218 186 219
rect 186 218 187 219
rect 187 218 188 219
rect 188 218 189 219
rect 189 218 190 219
rect 108 217 109 218
rect 109 217 110 218
rect 110 217 111 218
rect 111 217 112 218
rect 112 217 113 218
rect 113 217 114 218
rect 114 217 115 218
rect 115 217 116 218
rect 116 217 117 218
rect 117 217 118 218
rect 118 217 119 218
rect 119 217 120 218
rect 120 217 121 218
rect 121 217 122 218
rect 122 217 123 218
rect 123 217 124 218
rect 124 217 125 218
rect 125 217 126 218
rect 126 217 127 218
rect 127 217 128 218
rect 128 217 129 218
rect 168 217 169 218
rect 169 217 170 218
rect 170 217 171 218
rect 171 217 172 218
rect 172 217 173 218
rect 173 217 174 218
rect 174 217 175 218
rect 175 217 176 218
rect 176 217 177 218
rect 177 217 178 218
rect 178 217 179 218
rect 179 217 180 218
rect 180 217 181 218
rect 181 217 182 218
rect 182 217 183 218
rect 183 217 184 218
rect 184 217 185 218
rect 185 217 186 218
rect 186 217 187 218
rect 187 217 188 218
rect 188 217 189 218
rect 189 217 190 218
rect 104 216 105 217
rect 105 216 106 217
rect 106 216 107 217
rect 107 216 108 217
rect 108 216 109 217
rect 109 216 110 217
rect 110 216 111 217
rect 111 216 112 217
rect 112 216 113 217
rect 113 216 114 217
rect 114 216 115 217
rect 115 216 116 217
rect 116 216 117 217
rect 117 216 118 217
rect 118 216 119 217
rect 119 216 120 217
rect 120 216 121 217
rect 121 216 122 217
rect 122 216 123 217
rect 123 216 124 217
rect 124 216 125 217
rect 125 216 126 217
rect 126 216 127 217
rect 127 216 128 217
rect 128 216 129 217
rect 129 216 130 217
rect 130 216 131 217
rect 131 216 132 217
rect 132 216 133 217
rect 133 216 134 217
rect 134 216 135 217
rect 135 216 136 217
rect 136 216 137 217
rect 167 216 168 217
rect 168 216 169 217
rect 169 216 170 217
rect 170 216 171 217
rect 171 216 172 217
rect 172 216 173 217
rect 173 216 174 217
rect 174 216 175 217
rect 175 216 176 217
rect 176 216 177 217
rect 177 216 178 217
rect 178 216 179 217
rect 179 216 180 217
rect 180 216 181 217
rect 181 216 182 217
rect 182 216 183 217
rect 183 216 184 217
rect 184 216 185 217
rect 185 216 186 217
rect 186 216 187 217
rect 187 216 188 217
rect 188 216 189 217
rect 189 216 190 217
rect 103 215 104 216
rect 104 215 105 216
rect 105 215 106 216
rect 106 215 107 216
rect 107 215 108 216
rect 108 215 109 216
rect 109 215 110 216
rect 110 215 111 216
rect 111 215 112 216
rect 112 215 113 216
rect 113 215 114 216
rect 114 215 115 216
rect 115 215 116 216
rect 117 215 118 216
rect 118 215 119 216
rect 119 215 120 216
rect 120 215 121 216
rect 121 215 122 216
rect 124 215 125 216
rect 125 215 126 216
rect 126 215 127 216
rect 127 215 128 216
rect 128 215 129 216
rect 129 215 130 216
rect 130 215 131 216
rect 131 215 132 216
rect 132 215 133 216
rect 133 215 134 216
rect 134 215 135 216
rect 135 215 136 216
rect 136 215 137 216
rect 137 215 138 216
rect 138 215 139 216
rect 139 215 140 216
rect 166 215 167 216
rect 167 215 168 216
rect 168 215 169 216
rect 169 215 170 216
rect 170 215 171 216
rect 171 215 172 216
rect 172 215 173 216
rect 173 215 174 216
rect 174 215 175 216
rect 175 215 176 216
rect 176 215 177 216
rect 177 215 178 216
rect 178 215 179 216
rect 179 215 180 216
rect 180 215 181 216
rect 181 215 182 216
rect 182 215 183 216
rect 183 215 184 216
rect 184 215 185 216
rect 185 215 186 216
rect 186 215 187 216
rect 187 215 188 216
rect 188 215 189 216
rect 189 215 190 216
rect 101 214 102 215
rect 102 214 103 215
rect 103 214 104 215
rect 104 214 105 215
rect 105 214 106 215
rect 106 214 107 215
rect 107 214 108 215
rect 108 214 109 215
rect 109 214 110 215
rect 110 214 111 215
rect 111 214 112 215
rect 130 214 131 215
rect 131 214 132 215
rect 132 214 133 215
rect 133 214 134 215
rect 134 214 135 215
rect 135 214 136 215
rect 136 214 137 215
rect 137 214 138 215
rect 138 214 139 215
rect 139 214 140 215
rect 140 214 141 215
rect 165 214 166 215
rect 166 214 167 215
rect 167 214 168 215
rect 168 214 169 215
rect 169 214 170 215
rect 170 214 171 215
rect 171 214 172 215
rect 172 214 173 215
rect 173 214 174 215
rect 176 214 177 215
rect 177 214 178 215
rect 178 214 179 215
rect 179 214 180 215
rect 180 214 181 215
rect 181 214 182 215
rect 182 214 183 215
rect 183 214 184 215
rect 184 214 185 215
rect 185 214 186 215
rect 186 214 187 215
rect 187 214 188 215
rect 188 214 189 215
rect 189 214 190 215
rect 100 213 101 214
rect 101 213 102 214
rect 102 213 103 214
rect 103 213 104 214
rect 104 213 105 214
rect 105 213 106 214
rect 106 213 107 214
rect 133 213 134 214
rect 134 213 135 214
rect 135 213 136 214
rect 136 213 137 214
rect 137 213 138 214
rect 138 213 139 214
rect 139 213 140 214
rect 140 213 141 214
rect 141 213 142 214
rect 164 213 165 214
rect 165 213 166 214
rect 166 213 167 214
rect 167 213 168 214
rect 168 213 169 214
rect 169 213 170 214
rect 170 213 171 214
rect 171 213 172 214
rect 172 213 173 214
rect 176 213 177 214
rect 177 213 178 214
rect 178 213 179 214
rect 179 213 180 214
rect 180 213 181 214
rect 181 213 182 214
rect 182 213 183 214
rect 183 213 184 214
rect 184 213 185 214
rect 185 213 186 214
rect 186 213 187 214
rect 187 213 188 214
rect 188 213 189 214
rect 189 213 190 214
rect 99 212 100 213
rect 100 212 101 213
rect 101 212 102 213
rect 102 212 103 213
rect 103 212 104 213
rect 136 212 137 213
rect 137 212 138 213
rect 138 212 139 213
rect 139 212 140 213
rect 140 212 141 213
rect 141 212 142 213
rect 142 212 143 213
rect 143 212 144 213
rect 164 212 165 213
rect 165 212 166 213
rect 166 212 167 213
rect 167 212 168 213
rect 168 212 169 213
rect 169 212 170 213
rect 170 212 171 213
rect 171 212 172 213
rect 176 212 177 213
rect 177 212 178 213
rect 178 212 179 213
rect 179 212 180 213
rect 180 212 181 213
rect 181 212 182 213
rect 182 212 183 213
rect 183 212 184 213
rect 184 212 185 213
rect 185 212 186 213
rect 186 212 187 213
rect 187 212 188 213
rect 188 212 189 213
rect 189 212 190 213
rect 98 211 99 212
rect 99 211 100 212
rect 100 211 101 212
rect 101 211 102 212
rect 137 211 138 212
rect 138 211 139 212
rect 139 211 140 212
rect 140 211 141 212
rect 141 211 142 212
rect 142 211 143 212
rect 143 211 144 212
rect 144 211 145 212
rect 163 211 164 212
rect 164 211 165 212
rect 165 211 166 212
rect 166 211 167 212
rect 167 211 168 212
rect 168 211 169 212
rect 169 211 170 212
rect 170 211 171 212
rect 176 211 177 212
rect 177 211 178 212
rect 178 211 179 212
rect 179 211 180 212
rect 180 211 181 212
rect 181 211 182 212
rect 182 211 183 212
rect 183 211 184 212
rect 184 211 185 212
rect 185 211 186 212
rect 186 211 187 212
rect 187 211 188 212
rect 188 211 189 212
rect 189 211 190 212
rect 98 210 99 211
rect 99 210 100 211
rect 139 210 140 211
rect 140 210 141 211
rect 141 210 142 211
rect 142 210 143 211
rect 143 210 144 211
rect 144 210 145 211
rect 162 210 163 211
rect 163 210 164 211
rect 164 210 165 211
rect 165 210 166 211
rect 166 210 167 211
rect 167 210 168 211
rect 168 210 169 211
rect 169 210 170 211
rect 176 210 177 211
rect 177 210 178 211
rect 178 210 179 211
rect 179 210 180 211
rect 180 210 181 211
rect 181 210 182 211
rect 182 210 183 211
rect 183 210 184 211
rect 184 210 185 211
rect 185 210 186 211
rect 186 210 187 211
rect 187 210 188 211
rect 188 210 189 211
rect 189 210 190 211
rect 95 209 96 210
rect 140 209 141 210
rect 141 209 142 210
rect 142 209 143 210
rect 143 209 144 210
rect 144 209 145 210
rect 145 209 146 210
rect 146 209 147 210
rect 147 209 148 210
rect 160 209 161 210
rect 161 209 162 210
rect 162 209 163 210
rect 163 209 164 210
rect 164 209 165 210
rect 165 209 166 210
rect 166 209 167 210
rect 167 209 168 210
rect 168 209 169 210
rect 176 209 177 210
rect 177 209 178 210
rect 178 209 179 210
rect 179 209 180 210
rect 180 209 181 210
rect 181 209 182 210
rect 182 209 183 210
rect 183 209 184 210
rect 184 209 185 210
rect 185 209 186 210
rect 186 209 187 210
rect 187 209 188 210
rect 188 209 189 210
rect 189 209 190 210
rect 94 208 95 209
rect 95 208 96 209
rect 143 208 144 209
rect 144 208 145 209
rect 145 208 146 209
rect 146 208 147 209
rect 147 208 148 209
rect 148 208 149 209
rect 160 208 161 209
rect 161 208 162 209
rect 162 208 163 209
rect 163 208 164 209
rect 164 208 165 209
rect 165 208 166 209
rect 166 208 167 209
rect 176 208 177 209
rect 177 208 178 209
rect 178 208 179 209
rect 179 208 180 209
rect 180 208 181 209
rect 181 208 182 209
rect 182 208 183 209
rect 183 208 184 209
rect 184 208 185 209
rect 185 208 186 209
rect 186 208 187 209
rect 187 208 188 209
rect 188 208 189 209
rect 189 208 190 209
rect 93 207 94 208
rect 94 207 95 208
rect 95 207 96 208
rect 144 207 145 208
rect 145 207 146 208
rect 146 207 147 208
rect 147 207 148 208
rect 148 207 149 208
rect 159 207 160 208
rect 160 207 161 208
rect 161 207 162 208
rect 162 207 163 208
rect 163 207 164 208
rect 164 207 165 208
rect 165 207 166 208
rect 176 207 177 208
rect 177 207 178 208
rect 178 207 179 208
rect 179 207 180 208
rect 180 207 181 208
rect 181 207 182 208
rect 182 207 183 208
rect 183 207 184 208
rect 184 207 185 208
rect 185 207 186 208
rect 186 207 187 208
rect 187 207 188 208
rect 188 207 189 208
rect 189 207 190 208
rect 91 206 92 207
rect 92 206 93 207
rect 93 206 94 207
rect 94 206 95 207
rect 144 206 145 207
rect 145 206 146 207
rect 146 206 147 207
rect 147 206 148 207
rect 148 206 149 207
rect 149 206 150 207
rect 150 206 151 207
rect 158 206 159 207
rect 159 206 160 207
rect 160 206 161 207
rect 161 206 162 207
rect 162 206 163 207
rect 163 206 164 207
rect 164 206 165 207
rect 176 206 177 207
rect 177 206 178 207
rect 178 206 179 207
rect 179 206 180 207
rect 180 206 181 207
rect 181 206 182 207
rect 182 206 183 207
rect 183 206 184 207
rect 184 206 185 207
rect 185 206 186 207
rect 186 206 187 207
rect 187 206 188 207
rect 188 206 189 207
rect 189 206 190 207
rect 91 205 92 206
rect 92 205 93 206
rect 93 205 94 206
rect 145 205 146 206
rect 146 205 147 206
rect 147 205 148 206
rect 148 205 149 206
rect 149 205 150 206
rect 150 205 151 206
rect 151 205 152 206
rect 156 205 157 206
rect 157 205 158 206
rect 158 205 159 206
rect 159 205 160 206
rect 160 205 161 206
rect 161 205 162 206
rect 162 205 163 206
rect 163 205 164 206
rect 164 205 165 206
rect 176 205 177 206
rect 177 205 178 206
rect 178 205 179 206
rect 179 205 180 206
rect 180 205 181 206
rect 181 205 182 206
rect 182 205 183 206
rect 183 205 184 206
rect 184 205 185 206
rect 185 205 186 206
rect 186 205 187 206
rect 187 205 188 206
rect 188 205 189 206
rect 189 205 190 206
rect 91 204 92 205
rect 92 204 93 205
rect 146 204 147 205
rect 147 204 148 205
rect 148 204 149 205
rect 149 204 150 205
rect 150 204 151 205
rect 151 204 152 205
rect 152 204 153 205
rect 156 204 157 205
rect 157 204 158 205
rect 158 204 159 205
rect 159 204 160 205
rect 160 204 161 205
rect 161 204 162 205
rect 162 204 163 205
rect 163 204 164 205
rect 176 204 177 205
rect 177 204 178 205
rect 178 204 179 205
rect 179 204 180 205
rect 180 204 181 205
rect 181 204 182 205
rect 182 204 183 205
rect 183 204 184 205
rect 184 204 185 205
rect 185 204 186 205
rect 186 204 187 205
rect 187 204 188 205
rect 188 204 189 205
rect 90 203 91 204
rect 91 203 92 204
rect 147 203 148 204
rect 148 203 149 204
rect 149 203 150 204
rect 150 203 151 204
rect 151 203 152 204
rect 152 203 153 204
rect 153 203 154 204
rect 154 203 155 204
rect 155 203 156 204
rect 156 203 157 204
rect 157 203 158 204
rect 158 203 159 204
rect 159 203 160 204
rect 160 203 161 204
rect 161 203 162 204
rect 162 203 163 204
rect 176 203 177 204
rect 177 203 178 204
rect 178 203 179 204
rect 179 203 180 204
rect 180 203 181 204
rect 181 203 182 204
rect 182 203 183 204
rect 183 203 184 204
rect 184 203 185 204
rect 185 203 186 204
rect 186 203 187 204
rect 88 202 89 203
rect 89 202 90 203
rect 90 202 91 203
rect 91 202 92 203
rect 148 202 149 203
rect 149 202 150 203
rect 150 202 151 203
rect 151 202 152 203
rect 152 202 153 203
rect 153 202 154 203
rect 154 202 155 203
rect 155 202 156 203
rect 156 202 157 203
rect 157 202 158 203
rect 158 202 159 203
rect 159 202 160 203
rect 160 202 161 203
rect 161 202 162 203
rect 162 202 163 203
rect 175 202 176 203
rect 176 202 177 203
rect 177 202 178 203
rect 178 202 179 203
rect 179 202 180 203
rect 180 202 181 203
rect 181 202 182 203
rect 182 202 183 203
rect 183 202 184 203
rect 184 202 185 203
rect 87 201 88 202
rect 88 201 89 202
rect 89 201 90 202
rect 148 201 149 202
rect 149 201 150 202
rect 150 201 151 202
rect 151 201 152 202
rect 152 201 153 202
rect 153 201 154 202
rect 154 201 155 202
rect 155 201 156 202
rect 156 201 157 202
rect 157 201 158 202
rect 158 201 159 202
rect 159 201 160 202
rect 160 201 161 202
rect 175 201 176 202
rect 176 201 177 202
rect 177 201 178 202
rect 178 201 179 202
rect 179 201 180 202
rect 180 201 181 202
rect 181 201 182 202
rect 87 200 88 201
rect 88 200 89 201
rect 89 200 90 201
rect 148 200 149 201
rect 149 200 150 201
rect 150 200 151 201
rect 151 200 152 201
rect 152 200 153 201
rect 153 200 154 201
rect 154 200 155 201
rect 155 200 156 201
rect 156 200 157 201
rect 157 200 158 201
rect 158 200 159 201
rect 159 200 160 201
rect 160 200 161 201
rect 174 200 175 201
rect 175 200 176 201
rect 176 200 177 201
rect 177 200 178 201
rect 178 200 179 201
rect 179 200 180 201
rect 180 200 181 201
rect 85 199 86 200
rect 86 199 87 200
rect 87 199 88 200
rect 88 199 89 200
rect 148 199 149 200
rect 149 199 150 200
rect 150 199 151 200
rect 151 199 152 200
rect 152 199 153 200
rect 153 199 154 200
rect 154 199 155 200
rect 155 199 156 200
rect 156 199 157 200
rect 157 199 158 200
rect 158 199 159 200
rect 159 199 160 200
rect 160 199 161 200
rect 174 199 175 200
rect 175 199 176 200
rect 176 199 177 200
rect 177 199 178 200
rect 178 199 179 200
rect 85 198 86 199
rect 86 198 87 199
rect 87 198 88 199
rect 148 198 149 199
rect 149 198 150 199
rect 150 198 151 199
rect 151 198 152 199
rect 152 198 153 199
rect 153 198 154 199
rect 154 198 155 199
rect 155 198 156 199
rect 156 198 157 199
rect 157 198 158 199
rect 158 198 159 199
rect 159 198 160 199
rect 172 198 173 199
rect 173 198 174 199
rect 174 198 175 199
rect 175 198 176 199
rect 176 198 177 199
rect 177 198 178 199
rect 83 197 84 198
rect 84 197 85 198
rect 85 197 86 198
rect 86 197 87 198
rect 148 197 149 198
rect 149 197 150 198
rect 150 197 151 198
rect 151 197 152 198
rect 152 197 153 198
rect 153 197 154 198
rect 154 197 155 198
rect 155 197 156 198
rect 156 197 157 198
rect 157 197 158 198
rect 158 197 159 198
rect 172 197 173 198
rect 173 197 174 198
rect 174 197 175 198
rect 175 197 176 198
rect 176 197 177 198
rect 83 196 84 197
rect 84 196 85 197
rect 85 196 86 197
rect 86 196 87 197
rect 147 196 148 197
rect 148 196 149 197
rect 149 196 150 197
rect 150 196 151 197
rect 151 196 152 197
rect 152 196 153 197
rect 153 196 154 197
rect 154 196 155 197
rect 155 196 156 197
rect 156 196 157 197
rect 157 196 158 197
rect 158 196 159 197
rect 170 196 171 197
rect 171 196 172 197
rect 172 196 173 197
rect 173 196 174 197
rect 174 196 175 197
rect 175 196 176 197
rect 81 195 82 196
rect 82 195 83 196
rect 83 195 84 196
rect 147 195 148 196
rect 148 195 149 196
rect 149 195 150 196
rect 150 195 151 196
rect 151 195 152 196
rect 152 195 153 196
rect 153 195 154 196
rect 154 195 155 196
rect 155 195 156 196
rect 156 195 157 196
rect 168 195 169 196
rect 169 195 170 196
rect 170 195 171 196
rect 171 195 172 196
rect 172 195 173 196
rect 80 194 81 195
rect 81 194 82 195
rect 82 194 83 195
rect 83 194 84 195
rect 146 194 147 195
rect 147 194 148 195
rect 148 194 149 195
rect 149 194 150 195
rect 150 194 151 195
rect 151 194 152 195
rect 152 194 153 195
rect 153 194 154 195
rect 154 194 155 195
rect 155 194 156 195
rect 156 194 157 195
rect 168 194 169 195
rect 169 194 170 195
rect 170 194 171 195
rect 171 194 172 195
rect 172 194 173 195
rect 79 193 80 194
rect 80 193 81 194
rect 81 193 82 194
rect 82 193 83 194
rect 83 193 84 194
rect 146 193 147 194
rect 147 193 148 194
rect 148 193 149 194
rect 149 193 150 194
rect 150 193 151 194
rect 151 193 152 194
rect 152 193 153 194
rect 153 193 154 194
rect 154 193 155 194
rect 155 193 156 194
rect 156 193 157 194
rect 167 193 168 194
rect 168 193 169 194
rect 169 193 170 194
rect 170 193 171 194
rect 79 192 80 193
rect 80 192 81 193
rect 81 192 82 193
rect 146 192 147 193
rect 147 192 148 193
rect 148 192 149 193
rect 149 192 150 193
rect 150 192 151 193
rect 151 192 152 193
rect 152 192 153 193
rect 153 192 154 193
rect 154 192 155 193
rect 155 192 156 193
rect 165 192 166 193
rect 166 192 167 193
rect 167 192 168 193
rect 168 192 169 193
rect 169 192 170 193
rect 170 192 171 193
rect 78 191 79 192
rect 79 191 80 192
rect 80 191 81 192
rect 146 191 147 192
rect 147 191 148 192
rect 148 191 149 192
rect 149 191 150 192
rect 150 191 151 192
rect 151 191 152 192
rect 152 191 153 192
rect 153 191 154 192
rect 154 191 155 192
rect 155 191 156 192
rect 164 191 165 192
rect 165 191 166 192
rect 166 191 167 192
rect 167 191 168 192
rect 168 191 169 192
rect 77 190 78 191
rect 78 190 79 191
rect 79 190 80 191
rect 146 190 147 191
rect 147 190 148 191
rect 148 190 149 191
rect 149 190 150 191
rect 150 190 151 191
rect 151 190 152 191
rect 152 190 153 191
rect 153 190 154 191
rect 154 190 155 191
rect 163 190 164 191
rect 164 190 165 191
rect 165 190 166 191
rect 166 190 167 191
rect 167 190 168 191
rect 168 190 169 191
rect 75 189 76 190
rect 76 189 77 190
rect 77 189 78 190
rect 78 189 79 190
rect 79 189 80 190
rect 145 189 146 190
rect 146 189 147 190
rect 147 189 148 190
rect 148 189 149 190
rect 149 189 150 190
rect 150 189 151 190
rect 151 189 152 190
rect 152 189 153 190
rect 153 189 154 190
rect 154 189 155 190
rect 160 189 161 190
rect 161 189 162 190
rect 162 189 163 190
rect 163 189 164 190
rect 164 189 165 190
rect 165 189 166 190
rect 166 189 167 190
rect 167 189 168 190
rect 74 188 75 189
rect 75 188 76 189
rect 76 188 77 189
rect 145 188 146 189
rect 146 188 147 189
rect 147 188 148 189
rect 148 188 149 189
rect 149 188 150 189
rect 150 188 151 189
rect 151 188 152 189
rect 152 188 153 189
rect 153 188 154 189
rect 160 188 161 189
rect 161 188 162 189
rect 162 188 163 189
rect 163 188 164 189
rect 164 188 165 189
rect 165 188 166 189
rect 73 187 74 188
rect 74 187 75 188
rect 75 187 76 188
rect 146 187 147 188
rect 147 187 148 188
rect 148 187 149 188
rect 149 187 150 188
rect 150 187 151 188
rect 151 187 152 188
rect 152 187 153 188
rect 153 187 154 188
rect 159 187 160 188
rect 160 187 161 188
rect 161 187 162 188
rect 162 187 163 188
rect 163 187 164 188
rect 164 187 165 188
rect 165 187 166 188
rect 72 186 73 187
rect 73 186 74 187
rect 74 186 75 187
rect 75 186 76 187
rect 146 186 147 187
rect 147 186 148 187
rect 148 186 149 187
rect 149 186 150 187
rect 150 186 151 187
rect 151 186 152 187
rect 152 186 153 187
rect 158 186 159 187
rect 159 186 160 187
rect 160 186 161 187
rect 161 186 162 187
rect 162 186 163 187
rect 163 186 164 187
rect 164 186 165 187
rect 71 185 72 186
rect 72 185 73 186
rect 73 185 74 186
rect 146 185 147 186
rect 147 185 148 186
rect 148 185 149 186
rect 149 185 150 186
rect 150 185 151 186
rect 151 185 152 186
rect 152 185 153 186
rect 157 185 158 186
rect 158 185 159 186
rect 159 185 160 186
rect 160 185 161 186
rect 161 185 162 186
rect 162 185 163 186
rect 163 185 164 186
rect 164 185 165 186
rect 71 184 72 185
rect 72 184 73 185
rect 145 184 146 185
rect 146 184 147 185
rect 147 184 148 185
rect 148 184 149 185
rect 149 184 150 185
rect 150 184 151 185
rect 151 184 152 185
rect 152 184 153 185
rect 156 184 157 185
rect 157 184 158 185
rect 158 184 159 185
rect 159 184 160 185
rect 160 184 161 185
rect 161 184 162 185
rect 162 184 163 185
rect 163 184 164 185
rect 69 183 70 184
rect 70 183 71 184
rect 71 183 72 184
rect 145 183 146 184
rect 146 183 147 184
rect 147 183 148 184
rect 148 183 149 184
rect 149 183 150 184
rect 150 183 151 184
rect 151 183 152 184
rect 152 183 153 184
rect 156 183 157 184
rect 157 183 158 184
rect 158 183 159 184
rect 159 183 160 184
rect 160 183 161 184
rect 161 183 162 184
rect 162 183 163 184
rect 67 182 68 183
rect 68 182 69 183
rect 69 182 70 183
rect 70 182 71 183
rect 71 182 72 183
rect 95 182 96 183
rect 96 182 97 183
rect 97 182 98 183
rect 98 182 99 183
rect 99 182 100 183
rect 100 182 101 183
rect 101 182 102 183
rect 102 182 103 183
rect 103 182 104 183
rect 104 182 105 183
rect 105 182 106 183
rect 106 182 107 183
rect 107 182 108 183
rect 108 182 109 183
rect 109 182 110 183
rect 110 182 111 183
rect 145 182 146 183
rect 146 182 147 183
rect 147 182 148 183
rect 148 182 149 183
rect 149 182 150 183
rect 150 182 151 183
rect 151 182 152 183
rect 152 182 153 183
rect 154 182 155 183
rect 155 182 156 183
rect 156 182 157 183
rect 157 182 158 183
rect 158 182 159 183
rect 159 182 160 183
rect 160 182 161 183
rect 161 182 162 183
rect 66 181 67 182
rect 67 181 68 182
rect 68 181 69 182
rect 92 181 93 182
rect 93 181 94 182
rect 94 181 95 182
rect 95 181 96 182
rect 96 181 97 182
rect 97 181 98 182
rect 98 181 99 182
rect 99 181 100 182
rect 100 181 101 182
rect 101 181 102 182
rect 102 181 103 182
rect 103 181 104 182
rect 104 181 105 182
rect 105 181 106 182
rect 106 181 107 182
rect 107 181 108 182
rect 108 181 109 182
rect 109 181 110 182
rect 110 181 111 182
rect 111 181 112 182
rect 112 181 113 182
rect 113 181 114 182
rect 114 181 115 182
rect 146 181 147 182
rect 147 181 148 182
rect 148 181 149 182
rect 149 181 150 182
rect 150 181 151 182
rect 151 181 152 182
rect 154 181 155 182
rect 155 181 156 182
rect 156 181 157 182
rect 157 181 158 182
rect 158 181 159 182
rect 159 181 160 182
rect 160 181 161 182
rect 65 180 66 181
rect 66 180 67 181
rect 67 180 68 181
rect 90 180 91 181
rect 91 180 92 181
rect 92 180 93 181
rect 93 180 94 181
rect 94 180 95 181
rect 95 180 96 181
rect 96 180 97 181
rect 97 180 98 181
rect 98 180 99 181
rect 99 180 100 181
rect 100 180 101 181
rect 101 180 102 181
rect 102 180 103 181
rect 103 180 104 181
rect 104 180 105 181
rect 105 180 106 181
rect 106 180 107 181
rect 107 180 108 181
rect 108 180 109 181
rect 109 180 110 181
rect 110 180 111 181
rect 111 180 112 181
rect 112 180 113 181
rect 113 180 114 181
rect 114 180 115 181
rect 115 180 116 181
rect 116 180 117 181
rect 117 180 118 181
rect 146 180 147 181
rect 147 180 148 181
rect 148 180 149 181
rect 149 180 150 181
rect 150 180 151 181
rect 151 180 152 181
rect 154 180 155 181
rect 155 180 156 181
rect 156 180 157 181
rect 157 180 158 181
rect 158 180 159 181
rect 159 180 160 181
rect 160 180 161 181
rect 64 179 65 180
rect 65 179 66 180
rect 66 179 67 180
rect 90 179 91 180
rect 91 179 92 180
rect 92 179 93 180
rect 93 179 94 180
rect 94 179 95 180
rect 95 179 96 180
rect 96 179 97 180
rect 99 179 100 180
rect 100 179 101 180
rect 103 179 104 180
rect 104 179 105 180
rect 105 179 106 180
rect 106 179 107 180
rect 107 179 108 180
rect 108 179 109 180
rect 109 179 110 180
rect 110 179 111 180
rect 111 179 112 180
rect 112 179 113 180
rect 113 179 114 180
rect 114 179 115 180
rect 115 179 116 180
rect 116 179 117 180
rect 117 179 118 180
rect 118 179 119 180
rect 119 179 120 180
rect 120 179 121 180
rect 145 179 146 180
rect 146 179 147 180
rect 147 179 148 180
rect 148 179 149 180
rect 149 179 150 180
rect 150 179 151 180
rect 151 179 152 180
rect 153 179 154 180
rect 154 179 155 180
rect 155 179 156 180
rect 156 179 157 180
rect 157 179 158 180
rect 158 179 159 180
rect 159 179 160 180
rect 160 179 161 180
rect 63 178 64 179
rect 64 178 65 179
rect 65 178 66 179
rect 110 178 111 179
rect 111 178 112 179
rect 112 178 113 179
rect 113 178 114 179
rect 114 178 115 179
rect 115 178 116 179
rect 116 178 117 179
rect 117 178 118 179
rect 118 178 119 179
rect 119 178 120 179
rect 120 178 121 179
rect 121 178 122 179
rect 122 178 123 179
rect 145 178 146 179
rect 146 178 147 179
rect 147 178 148 179
rect 148 178 149 179
rect 149 178 150 179
rect 150 178 151 179
rect 151 178 152 179
rect 152 178 153 179
rect 153 178 154 179
rect 154 178 155 179
rect 155 178 156 179
rect 156 178 157 179
rect 157 178 158 179
rect 158 178 159 179
rect 159 178 160 179
rect 61 177 62 178
rect 62 177 63 178
rect 63 177 64 178
rect 64 177 65 178
rect 85 177 86 178
rect 86 177 87 178
rect 114 177 115 178
rect 115 177 116 178
rect 116 177 117 178
rect 117 177 118 178
rect 118 177 119 178
rect 119 177 120 178
rect 120 177 121 178
rect 121 177 122 178
rect 122 177 123 178
rect 123 177 124 178
rect 124 177 125 178
rect 146 177 147 178
rect 147 177 148 178
rect 148 177 149 178
rect 149 177 150 178
rect 150 177 151 178
rect 152 177 153 178
rect 153 177 154 178
rect 154 177 155 178
rect 155 177 156 178
rect 156 177 157 178
rect 157 177 158 178
rect 158 177 159 178
rect 60 176 61 177
rect 61 176 62 177
rect 62 176 63 177
rect 63 176 64 177
rect 83 176 84 177
rect 84 176 85 177
rect 85 176 86 177
rect 86 176 87 177
rect 117 176 118 177
rect 118 176 119 177
rect 119 176 120 177
rect 120 176 121 177
rect 121 176 122 177
rect 122 176 123 177
rect 123 176 124 177
rect 124 176 125 177
rect 125 176 126 177
rect 126 176 127 177
rect 127 176 128 177
rect 145 176 146 177
rect 146 176 147 177
rect 147 176 148 177
rect 148 176 149 177
rect 149 176 150 177
rect 150 176 151 177
rect 152 176 153 177
rect 153 176 154 177
rect 154 176 155 177
rect 155 176 156 177
rect 156 176 157 177
rect 157 176 158 177
rect 158 176 159 177
rect 58 175 59 176
rect 59 175 60 176
rect 60 175 61 176
rect 61 175 62 176
rect 62 175 63 176
rect 80 175 81 176
rect 81 175 82 176
rect 82 175 83 176
rect 83 175 84 176
rect 84 175 85 176
rect 85 175 86 176
rect 120 175 121 176
rect 121 175 122 176
rect 122 175 123 176
rect 123 175 124 176
rect 124 175 125 176
rect 125 175 126 176
rect 126 175 127 176
rect 127 175 128 176
rect 128 175 129 176
rect 129 175 130 176
rect 130 175 131 176
rect 131 175 132 176
rect 145 175 146 176
rect 146 175 147 176
rect 147 175 148 176
rect 148 175 149 176
rect 149 175 150 176
rect 150 175 151 176
rect 152 175 153 176
rect 153 175 154 176
rect 154 175 155 176
rect 155 175 156 176
rect 156 175 157 176
rect 157 175 158 176
rect 56 174 57 175
rect 57 174 58 175
rect 58 174 59 175
rect 59 174 60 175
rect 60 174 61 175
rect 79 174 80 175
rect 80 174 81 175
rect 81 174 82 175
rect 82 174 83 175
rect 83 174 84 175
rect 84 174 85 175
rect 127 174 128 175
rect 128 174 129 175
rect 129 174 130 175
rect 130 174 131 175
rect 131 174 132 175
rect 132 174 133 175
rect 133 174 134 175
rect 146 174 147 175
rect 147 174 148 175
rect 148 174 149 175
rect 149 174 150 175
rect 150 174 151 175
rect 152 174 153 175
rect 153 174 154 175
rect 154 174 155 175
rect 155 174 156 175
rect 156 174 157 175
rect 157 174 158 175
rect 54 173 55 174
rect 55 173 56 174
rect 56 173 57 174
rect 57 173 58 174
rect 58 173 59 174
rect 78 173 79 174
rect 79 173 80 174
rect 80 173 81 174
rect 81 173 82 174
rect 82 173 83 174
rect 83 173 84 174
rect 129 173 130 174
rect 130 173 131 174
rect 131 173 132 174
rect 132 173 133 174
rect 133 173 134 174
rect 134 173 135 174
rect 135 173 136 174
rect 136 173 137 174
rect 145 173 146 174
rect 146 173 147 174
rect 147 173 148 174
rect 148 173 149 174
rect 149 173 150 174
rect 150 173 151 174
rect 152 173 153 174
rect 153 173 154 174
rect 154 173 155 174
rect 155 173 156 174
rect 156 173 157 174
rect 157 173 158 174
rect 53 172 54 173
rect 54 172 55 173
rect 55 172 56 173
rect 56 172 57 173
rect 57 172 58 173
rect 58 172 59 173
rect 77 172 78 173
rect 78 172 79 173
rect 79 172 80 173
rect 80 172 81 173
rect 81 172 82 173
rect 82 172 83 173
rect 83 172 84 173
rect 132 172 133 173
rect 133 172 134 173
rect 134 172 135 173
rect 135 172 136 173
rect 136 172 137 173
rect 137 172 138 173
rect 145 172 146 173
rect 146 172 147 173
rect 147 172 148 173
rect 148 172 149 173
rect 149 172 150 173
rect 150 172 151 173
rect 152 172 153 173
rect 153 172 154 173
rect 154 172 155 173
rect 155 172 156 173
rect 156 172 157 173
rect 157 172 158 173
rect 52 171 53 172
rect 53 171 54 172
rect 54 171 55 172
rect 55 171 56 172
rect 56 171 57 172
rect 75 171 76 172
rect 76 171 77 172
rect 77 171 78 172
rect 78 171 79 172
rect 79 171 80 172
rect 80 171 81 172
rect 81 171 82 172
rect 82 171 83 172
rect 135 171 136 172
rect 136 171 137 172
rect 137 171 138 172
rect 138 171 139 172
rect 139 171 140 172
rect 145 171 146 172
rect 146 171 147 172
rect 147 171 148 172
rect 148 171 149 172
rect 149 171 150 172
rect 150 171 151 172
rect 152 171 153 172
rect 153 171 154 172
rect 154 171 155 172
rect 155 171 156 172
rect 156 171 157 172
rect 157 171 158 172
rect 168 171 169 172
rect 169 171 170 172
rect 190 171 191 172
rect 191 171 192 172
rect 193 171 194 172
rect 194 171 195 172
rect 196 171 197 172
rect 197 171 198 172
rect 50 170 51 171
rect 51 170 52 171
rect 52 170 53 171
rect 53 170 54 171
rect 54 170 55 171
rect 55 170 56 171
rect 75 170 76 171
rect 76 170 77 171
rect 77 170 78 171
rect 78 170 79 171
rect 79 170 80 171
rect 80 170 81 171
rect 81 170 82 171
rect 138 170 139 171
rect 139 170 140 171
rect 145 170 146 171
rect 146 170 147 171
rect 147 170 148 171
rect 148 170 149 171
rect 149 170 150 171
rect 150 170 151 171
rect 152 170 153 171
rect 153 170 154 171
rect 154 170 155 171
rect 155 170 156 171
rect 156 170 157 171
rect 157 170 158 171
rect 165 170 166 171
rect 166 170 167 171
rect 167 170 168 171
rect 168 170 169 171
rect 169 170 170 171
rect 170 170 171 171
rect 171 170 172 171
rect 172 170 173 171
rect 173 170 174 171
rect 174 170 175 171
rect 175 170 176 171
rect 176 170 177 171
rect 177 170 178 171
rect 178 170 179 171
rect 179 170 180 171
rect 180 170 181 171
rect 181 170 182 171
rect 182 170 183 171
rect 183 170 184 171
rect 184 170 185 171
rect 185 170 186 171
rect 186 170 187 171
rect 187 170 188 171
rect 188 170 189 171
rect 189 170 190 171
rect 190 170 191 171
rect 191 170 192 171
rect 192 170 193 171
rect 193 170 194 171
rect 194 170 195 171
rect 195 170 196 171
rect 196 170 197 171
rect 197 170 198 171
rect 198 170 199 171
rect 199 170 200 171
rect 200 170 201 171
rect 201 170 202 171
rect 202 170 203 171
rect 203 170 204 171
rect 204 170 205 171
rect 205 170 206 171
rect 49 169 50 170
rect 50 169 51 170
rect 51 169 52 170
rect 52 169 53 170
rect 53 169 54 170
rect 54 169 55 170
rect 74 169 75 170
rect 75 169 76 170
rect 76 169 77 170
rect 77 169 78 170
rect 78 169 79 170
rect 79 169 80 170
rect 80 169 81 170
rect 146 169 147 170
rect 147 169 148 170
rect 148 169 149 170
rect 149 169 150 170
rect 150 169 151 170
rect 151 169 152 170
rect 152 169 153 170
rect 153 169 154 170
rect 154 169 155 170
rect 155 169 156 170
rect 156 169 157 170
rect 157 169 158 170
rect 164 169 165 170
rect 165 169 166 170
rect 166 169 167 170
rect 167 169 168 170
rect 168 169 169 170
rect 169 169 170 170
rect 170 169 171 170
rect 171 169 172 170
rect 172 169 173 170
rect 173 169 174 170
rect 174 169 175 170
rect 175 169 176 170
rect 176 169 177 170
rect 177 169 178 170
rect 178 169 179 170
rect 179 169 180 170
rect 180 169 181 170
rect 181 169 182 170
rect 182 169 183 170
rect 183 169 184 170
rect 184 169 185 170
rect 185 169 186 170
rect 186 169 187 170
rect 187 169 188 170
rect 188 169 189 170
rect 189 169 190 170
rect 190 169 191 170
rect 191 169 192 170
rect 192 169 193 170
rect 193 169 194 170
rect 194 169 195 170
rect 195 169 196 170
rect 196 169 197 170
rect 197 169 198 170
rect 198 169 199 170
rect 199 169 200 170
rect 200 169 201 170
rect 201 169 202 170
rect 202 169 203 170
rect 203 169 204 170
rect 204 169 205 170
rect 205 169 206 170
rect 206 169 207 170
rect 207 169 208 170
rect 208 169 209 170
rect 209 169 210 170
rect 46 168 47 169
rect 47 168 48 169
rect 48 168 49 169
rect 49 168 50 169
rect 50 168 51 169
rect 51 168 52 169
rect 52 168 53 169
rect 53 168 54 169
rect 71 168 72 169
rect 72 168 73 169
rect 73 168 74 169
rect 74 168 75 169
rect 75 168 76 169
rect 76 168 77 169
rect 77 168 78 169
rect 78 168 79 169
rect 79 168 80 169
rect 145 168 146 169
rect 146 168 147 169
rect 147 168 148 169
rect 148 168 149 169
rect 149 168 150 169
rect 150 168 151 169
rect 151 168 152 169
rect 152 168 153 169
rect 153 168 154 169
rect 154 168 155 169
rect 155 168 156 169
rect 156 168 157 169
rect 157 168 158 169
rect 162 168 163 169
rect 163 168 164 169
rect 164 168 165 169
rect 165 168 166 169
rect 166 168 167 169
rect 167 168 168 169
rect 168 168 169 169
rect 169 168 170 169
rect 170 168 171 169
rect 171 168 172 169
rect 172 168 173 169
rect 173 168 174 169
rect 174 168 175 169
rect 175 168 176 169
rect 176 168 177 169
rect 177 168 178 169
rect 178 168 179 169
rect 179 168 180 169
rect 180 168 181 169
rect 181 168 182 169
rect 182 168 183 169
rect 183 168 184 169
rect 184 168 185 169
rect 185 168 186 169
rect 186 168 187 169
rect 187 168 188 169
rect 188 168 189 169
rect 189 168 190 169
rect 190 168 191 169
rect 191 168 192 169
rect 192 168 193 169
rect 193 168 194 169
rect 194 168 195 169
rect 195 168 196 169
rect 196 168 197 169
rect 197 168 198 169
rect 198 168 199 169
rect 199 168 200 169
rect 200 168 201 169
rect 201 168 202 169
rect 202 168 203 169
rect 203 168 204 169
rect 204 168 205 169
rect 205 168 206 169
rect 206 168 207 169
rect 207 168 208 169
rect 208 168 209 169
rect 209 168 210 169
rect 210 168 211 169
rect 211 168 212 169
rect 212 168 213 169
rect 213 168 214 169
rect 44 167 45 168
rect 45 167 46 168
rect 46 167 47 168
rect 47 167 48 168
rect 48 167 49 168
rect 49 167 50 168
rect 50 167 51 168
rect 51 167 52 168
rect 71 167 72 168
rect 72 167 73 168
rect 73 167 74 168
rect 74 167 75 168
rect 75 167 76 168
rect 76 167 77 168
rect 77 167 78 168
rect 78 167 79 168
rect 145 167 146 168
rect 146 167 147 168
rect 147 167 148 168
rect 148 167 149 168
rect 149 167 150 168
rect 150 167 151 168
rect 151 167 152 168
rect 152 167 153 168
rect 153 167 154 168
rect 154 167 155 168
rect 155 167 156 168
rect 156 167 157 168
rect 157 167 158 168
rect 161 167 162 168
rect 162 167 163 168
rect 163 167 164 168
rect 164 167 165 168
rect 165 167 166 168
rect 166 167 167 168
rect 167 167 168 168
rect 168 167 169 168
rect 169 167 170 168
rect 170 167 171 168
rect 171 167 172 168
rect 172 167 173 168
rect 173 167 174 168
rect 174 167 175 168
rect 175 167 176 168
rect 176 167 177 168
rect 177 167 178 168
rect 178 167 179 168
rect 179 167 180 168
rect 180 167 181 168
rect 181 167 182 168
rect 182 167 183 168
rect 183 167 184 168
rect 199 167 200 168
rect 200 167 201 168
rect 201 167 202 168
rect 202 167 203 168
rect 203 167 204 168
rect 204 167 205 168
rect 205 167 206 168
rect 206 167 207 168
rect 207 167 208 168
rect 208 167 209 168
rect 209 167 210 168
rect 210 167 211 168
rect 211 167 212 168
rect 212 167 213 168
rect 213 167 214 168
rect 214 167 215 168
rect 215 167 216 168
rect 42 166 43 167
rect 43 166 44 167
rect 44 166 45 167
rect 45 166 46 167
rect 46 166 47 167
rect 47 166 48 167
rect 48 166 49 167
rect 49 166 50 167
rect 50 166 51 167
rect 70 166 71 167
rect 71 166 72 167
rect 72 166 73 167
rect 73 166 74 167
rect 74 166 75 167
rect 75 166 76 167
rect 76 166 77 167
rect 77 166 78 167
rect 145 166 146 167
rect 146 166 147 167
rect 147 166 148 167
rect 148 166 149 167
rect 149 166 150 167
rect 150 166 151 167
rect 151 166 152 167
rect 152 166 153 167
rect 153 166 154 167
rect 154 166 155 167
rect 155 166 156 167
rect 156 166 157 167
rect 157 166 158 167
rect 160 166 161 167
rect 161 166 162 167
rect 162 166 163 167
rect 163 166 164 167
rect 164 166 165 167
rect 165 166 166 167
rect 166 166 167 167
rect 167 166 168 167
rect 168 166 169 167
rect 169 166 170 167
rect 170 166 171 167
rect 171 166 172 167
rect 172 166 173 167
rect 173 166 174 167
rect 174 166 175 167
rect 175 166 176 167
rect 176 166 177 167
rect 177 166 178 167
rect 178 166 179 167
rect 179 166 180 167
rect 201 166 202 167
rect 202 166 203 167
rect 203 166 204 167
rect 204 166 205 167
rect 205 166 206 167
rect 206 166 207 167
rect 207 166 208 167
rect 208 166 209 167
rect 209 166 210 167
rect 210 166 211 167
rect 211 166 212 167
rect 212 166 213 167
rect 213 166 214 167
rect 214 166 215 167
rect 215 166 216 167
rect 216 166 217 167
rect 217 166 218 167
rect 42 165 43 166
rect 43 165 44 166
rect 44 165 45 166
rect 45 165 46 166
rect 46 165 47 166
rect 47 165 48 166
rect 48 165 49 166
rect 69 165 70 166
rect 70 165 71 166
rect 71 165 72 166
rect 72 165 73 166
rect 73 165 74 166
rect 74 165 75 166
rect 75 165 76 166
rect 76 165 77 166
rect 145 165 146 166
rect 146 165 147 166
rect 147 165 148 166
rect 148 165 149 166
rect 149 165 150 166
rect 150 165 151 166
rect 151 165 152 166
rect 152 165 153 166
rect 153 165 154 166
rect 154 165 155 166
rect 155 165 156 166
rect 156 165 157 166
rect 157 165 158 166
rect 158 165 159 166
rect 159 165 160 166
rect 160 165 161 166
rect 161 165 162 166
rect 162 165 163 166
rect 163 165 164 166
rect 164 165 165 166
rect 165 165 166 166
rect 166 165 167 166
rect 167 165 168 166
rect 168 165 169 166
rect 169 165 170 166
rect 170 165 171 166
rect 171 165 172 166
rect 172 165 173 166
rect 173 165 174 166
rect 174 165 175 166
rect 175 165 176 166
rect 176 165 177 166
rect 203 165 204 166
rect 204 165 205 166
rect 205 165 206 166
rect 206 165 207 166
rect 207 165 208 166
rect 208 165 209 166
rect 209 165 210 166
rect 210 165 211 166
rect 211 165 212 166
rect 212 165 213 166
rect 213 165 214 166
rect 214 165 215 166
rect 215 165 216 166
rect 216 165 217 166
rect 217 165 218 166
rect 39 164 40 165
rect 40 164 41 165
rect 41 164 42 165
rect 42 164 43 165
rect 43 164 44 165
rect 44 164 45 165
rect 45 164 46 165
rect 46 164 47 165
rect 47 164 48 165
rect 67 164 68 165
rect 68 164 69 165
rect 69 164 70 165
rect 70 164 71 165
rect 71 164 72 165
rect 72 164 73 165
rect 73 164 74 165
rect 74 164 75 165
rect 75 164 76 165
rect 145 164 146 165
rect 146 164 147 165
rect 147 164 148 165
rect 148 164 149 165
rect 149 164 150 165
rect 150 164 151 165
rect 151 164 152 165
rect 152 164 153 165
rect 153 164 154 165
rect 154 164 155 165
rect 155 164 156 165
rect 156 164 157 165
rect 157 164 158 165
rect 158 164 159 165
rect 159 164 160 165
rect 160 164 161 165
rect 161 164 162 165
rect 162 164 163 165
rect 163 164 164 165
rect 164 164 165 165
rect 165 164 166 165
rect 166 164 167 165
rect 167 164 168 165
rect 168 164 169 165
rect 169 164 170 165
rect 170 164 171 165
rect 171 164 172 165
rect 172 164 173 165
rect 173 164 174 165
rect 204 164 205 165
rect 205 164 206 165
rect 206 164 207 165
rect 207 164 208 165
rect 208 164 209 165
rect 209 164 210 165
rect 210 164 211 165
rect 211 164 212 165
rect 212 164 213 165
rect 213 164 214 165
rect 214 164 215 165
rect 215 164 216 165
rect 216 164 217 165
rect 217 164 218 165
rect 218 164 219 165
rect 219 164 220 165
rect 38 163 39 164
rect 39 163 40 164
rect 40 163 41 164
rect 41 163 42 164
rect 42 163 43 164
rect 43 163 44 164
rect 44 163 45 164
rect 45 163 46 164
rect 46 163 47 164
rect 67 163 68 164
rect 68 163 69 164
rect 69 163 70 164
rect 70 163 71 164
rect 71 163 72 164
rect 72 163 73 164
rect 73 163 74 164
rect 74 163 75 164
rect 75 163 76 164
rect 144 163 145 164
rect 145 163 146 164
rect 146 163 147 164
rect 147 163 148 164
rect 148 163 149 164
rect 149 163 150 164
rect 150 163 151 164
rect 151 163 152 164
rect 152 163 153 164
rect 153 163 154 164
rect 154 163 155 164
rect 155 163 156 164
rect 156 163 157 164
rect 157 163 158 164
rect 158 163 159 164
rect 159 163 160 164
rect 160 163 161 164
rect 161 163 162 164
rect 162 163 163 164
rect 163 163 164 164
rect 164 163 165 164
rect 165 163 166 164
rect 166 163 167 164
rect 167 163 168 164
rect 168 163 169 164
rect 169 163 170 164
rect 170 163 171 164
rect 205 163 206 164
rect 206 163 207 164
rect 207 163 208 164
rect 208 163 209 164
rect 209 163 210 164
rect 210 163 211 164
rect 211 163 212 164
rect 212 163 213 164
rect 213 163 214 164
rect 214 163 215 164
rect 215 163 216 164
rect 216 163 217 164
rect 217 163 218 164
rect 218 163 219 164
rect 219 163 220 164
rect 220 163 221 164
rect 36 162 37 163
rect 37 162 38 163
rect 38 162 39 163
rect 39 162 40 163
rect 40 162 41 163
rect 41 162 42 163
rect 42 162 43 163
rect 43 162 44 163
rect 44 162 45 163
rect 45 162 46 163
rect 66 162 67 163
rect 67 162 68 163
rect 68 162 69 163
rect 69 162 70 163
rect 70 162 71 163
rect 71 162 72 163
rect 72 162 73 163
rect 73 162 74 163
rect 74 162 75 163
rect 144 162 145 163
rect 145 162 146 163
rect 146 162 147 163
rect 147 162 148 163
rect 148 162 149 163
rect 149 162 150 163
rect 150 162 151 163
rect 151 162 152 163
rect 152 162 153 163
rect 153 162 154 163
rect 154 162 155 163
rect 155 162 156 163
rect 156 162 157 163
rect 157 162 158 163
rect 158 162 159 163
rect 159 162 160 163
rect 160 162 161 163
rect 161 162 162 163
rect 162 162 163 163
rect 163 162 164 163
rect 164 162 165 163
rect 165 162 166 163
rect 166 162 167 163
rect 167 162 168 163
rect 168 162 169 163
rect 206 162 207 163
rect 207 162 208 163
rect 208 162 209 163
rect 209 162 210 163
rect 210 162 211 163
rect 211 162 212 163
rect 212 162 213 163
rect 213 162 214 163
rect 214 162 215 163
rect 215 162 216 163
rect 216 162 217 163
rect 217 162 218 163
rect 218 162 219 163
rect 219 162 220 163
rect 220 162 221 163
rect 221 162 222 163
rect 33 161 34 162
rect 34 161 35 162
rect 35 161 36 162
rect 36 161 37 162
rect 37 161 38 162
rect 38 161 39 162
rect 39 161 40 162
rect 40 161 41 162
rect 41 161 42 162
rect 42 161 43 162
rect 43 161 44 162
rect 64 161 65 162
rect 65 161 66 162
rect 66 161 67 162
rect 67 161 68 162
rect 68 161 69 162
rect 69 161 70 162
rect 70 161 71 162
rect 71 161 72 162
rect 72 161 73 162
rect 73 161 74 162
rect 144 161 145 162
rect 145 161 146 162
rect 146 161 147 162
rect 147 161 148 162
rect 148 161 149 162
rect 149 161 150 162
rect 150 161 151 162
rect 151 161 152 162
rect 152 161 153 162
rect 153 161 154 162
rect 154 161 155 162
rect 155 161 156 162
rect 156 161 157 162
rect 157 161 158 162
rect 158 161 159 162
rect 159 161 160 162
rect 160 161 161 162
rect 161 161 162 162
rect 162 161 163 162
rect 163 161 164 162
rect 164 161 165 162
rect 208 161 209 162
rect 209 161 210 162
rect 210 161 211 162
rect 211 161 212 162
rect 212 161 213 162
rect 213 161 214 162
rect 214 161 215 162
rect 215 161 216 162
rect 216 161 217 162
rect 217 161 218 162
rect 218 161 219 162
rect 219 161 220 162
rect 220 161 221 162
rect 221 161 222 162
rect 222 161 223 162
rect 31 160 32 161
rect 32 160 33 161
rect 33 160 34 161
rect 34 160 35 161
rect 35 160 36 161
rect 36 160 37 161
rect 37 160 38 161
rect 38 160 39 161
rect 39 160 40 161
rect 40 160 41 161
rect 63 160 64 161
rect 64 160 65 161
rect 65 160 66 161
rect 66 160 67 161
rect 67 160 68 161
rect 68 160 69 161
rect 69 160 70 161
rect 70 160 71 161
rect 71 160 72 161
rect 143 160 144 161
rect 144 160 145 161
rect 145 160 146 161
rect 146 160 147 161
rect 147 160 148 161
rect 148 160 149 161
rect 149 160 150 161
rect 150 160 151 161
rect 151 160 152 161
rect 152 160 153 161
rect 153 160 154 161
rect 154 160 155 161
rect 155 160 156 161
rect 156 160 157 161
rect 157 160 158 161
rect 158 160 159 161
rect 159 160 160 161
rect 209 160 210 161
rect 210 160 211 161
rect 211 160 212 161
rect 212 160 213 161
rect 213 160 214 161
rect 214 160 215 161
rect 215 160 216 161
rect 216 160 217 161
rect 217 160 218 161
rect 218 160 219 161
rect 219 160 220 161
rect 220 160 221 161
rect 221 160 222 161
rect 222 160 223 161
rect 223 160 224 161
rect 29 159 30 160
rect 30 159 31 160
rect 31 159 32 160
rect 32 159 33 160
rect 33 159 34 160
rect 34 159 35 160
rect 35 159 36 160
rect 36 159 37 160
rect 37 159 38 160
rect 38 159 39 160
rect 63 159 64 160
rect 64 159 65 160
rect 65 159 66 160
rect 66 159 67 160
rect 67 159 68 160
rect 68 159 69 160
rect 69 159 70 160
rect 70 159 71 160
rect 71 159 72 160
rect 143 159 144 160
rect 144 159 145 160
rect 145 159 146 160
rect 146 159 147 160
rect 147 159 148 160
rect 148 159 149 160
rect 149 159 150 160
rect 150 159 151 160
rect 151 159 152 160
rect 152 159 153 160
rect 153 159 154 160
rect 154 159 155 160
rect 155 159 156 160
rect 156 159 157 160
rect 210 159 211 160
rect 211 159 212 160
rect 212 159 213 160
rect 213 159 214 160
rect 214 159 215 160
rect 215 159 216 160
rect 216 159 217 160
rect 217 159 218 160
rect 218 159 219 160
rect 219 159 220 160
rect 220 159 221 160
rect 221 159 222 160
rect 222 159 223 160
rect 223 159 224 160
rect 28 158 29 159
rect 29 158 30 159
rect 30 158 31 159
rect 31 158 32 159
rect 32 158 33 159
rect 33 158 34 159
rect 34 158 35 159
rect 35 158 36 159
rect 36 158 37 159
rect 37 158 38 159
rect 62 158 63 159
rect 63 158 64 159
rect 64 158 65 159
rect 65 158 66 159
rect 66 158 67 159
rect 67 158 68 159
rect 68 158 69 159
rect 69 158 70 159
rect 70 158 71 159
rect 142 158 143 159
rect 143 158 144 159
rect 144 158 145 159
rect 145 158 146 159
rect 146 158 147 159
rect 147 158 148 159
rect 148 158 149 159
rect 149 158 150 159
rect 150 158 151 159
rect 151 158 152 159
rect 152 158 153 159
rect 211 158 212 159
rect 212 158 213 159
rect 213 158 214 159
rect 214 158 215 159
rect 215 158 216 159
rect 216 158 217 159
rect 217 158 218 159
rect 218 158 219 159
rect 219 158 220 159
rect 220 158 221 159
rect 221 158 222 159
rect 222 158 223 159
rect 223 158 224 159
rect 224 158 225 159
rect 26 157 27 158
rect 27 157 28 158
rect 28 157 29 158
rect 29 157 30 158
rect 30 157 31 158
rect 31 157 32 158
rect 32 157 33 158
rect 33 157 34 158
rect 34 157 35 158
rect 35 157 36 158
rect 36 157 37 158
rect 61 157 62 158
rect 62 157 63 158
rect 63 157 64 158
rect 64 157 65 158
rect 65 157 66 158
rect 66 157 67 158
rect 67 157 68 158
rect 68 157 69 158
rect 141 157 142 158
rect 142 157 143 158
rect 143 157 144 158
rect 144 157 145 158
rect 145 157 146 158
rect 146 157 147 158
rect 147 157 148 158
rect 148 157 149 158
rect 212 157 213 158
rect 213 157 214 158
rect 214 157 215 158
rect 215 157 216 158
rect 216 157 217 158
rect 217 157 218 158
rect 218 157 219 158
rect 219 157 220 158
rect 220 157 221 158
rect 221 157 222 158
rect 222 157 223 158
rect 223 157 224 158
rect 224 157 225 158
rect 225 157 226 158
rect 24 156 25 157
rect 25 156 26 157
rect 26 156 27 157
rect 27 156 28 157
rect 28 156 29 157
rect 29 156 30 157
rect 30 156 31 157
rect 31 156 32 157
rect 32 156 33 157
rect 33 156 34 157
rect 34 156 35 157
rect 60 156 61 157
rect 61 156 62 157
rect 62 156 63 157
rect 63 156 64 157
rect 64 156 65 157
rect 65 156 66 157
rect 66 156 67 157
rect 67 156 68 157
rect 68 156 69 157
rect 141 156 142 157
rect 142 156 143 157
rect 144 156 145 157
rect 213 156 214 157
rect 214 156 215 157
rect 215 156 216 157
rect 216 156 217 157
rect 217 156 218 157
rect 218 156 219 157
rect 219 156 220 157
rect 220 156 221 157
rect 221 156 222 157
rect 222 156 223 157
rect 223 156 224 157
rect 224 156 225 157
rect 225 156 226 157
rect 20 155 21 156
rect 21 155 22 156
rect 22 155 23 156
rect 23 155 24 156
rect 24 155 25 156
rect 25 155 26 156
rect 26 155 27 156
rect 27 155 28 156
rect 28 155 29 156
rect 29 155 30 156
rect 30 155 31 156
rect 31 155 32 156
rect 32 155 33 156
rect 58 155 59 156
rect 59 155 60 156
rect 60 155 61 156
rect 61 155 62 156
rect 62 155 63 156
rect 63 155 64 156
rect 64 155 65 156
rect 65 155 66 156
rect 66 155 67 156
rect 67 155 68 156
rect 213 155 214 156
rect 214 155 215 156
rect 215 155 216 156
rect 216 155 217 156
rect 217 155 218 156
rect 218 155 219 156
rect 219 155 220 156
rect 220 155 221 156
rect 221 155 222 156
rect 222 155 223 156
rect 223 155 224 156
rect 224 155 225 156
rect 225 155 226 156
rect 18 154 19 155
rect 19 154 20 155
rect 20 154 21 155
rect 21 154 22 155
rect 22 154 23 155
rect 23 154 24 155
rect 24 154 25 155
rect 25 154 26 155
rect 26 154 27 155
rect 27 154 28 155
rect 28 154 29 155
rect 29 154 30 155
rect 58 154 59 155
rect 59 154 60 155
rect 60 154 61 155
rect 61 154 62 155
rect 62 154 63 155
rect 63 154 64 155
rect 64 154 65 155
rect 65 154 66 155
rect 66 154 67 155
rect 214 154 215 155
rect 215 154 216 155
rect 216 154 217 155
rect 217 154 218 155
rect 218 154 219 155
rect 219 154 220 155
rect 220 154 221 155
rect 221 154 222 155
rect 222 154 223 155
rect 223 154 224 155
rect 224 154 225 155
rect 225 154 226 155
rect 226 154 227 155
rect 17 153 18 154
rect 18 153 19 154
rect 19 153 20 154
rect 20 153 21 154
rect 21 153 22 154
rect 22 153 23 154
rect 23 153 24 154
rect 24 153 25 154
rect 25 153 26 154
rect 26 153 27 154
rect 57 153 58 154
rect 58 153 59 154
rect 59 153 60 154
rect 60 153 61 154
rect 61 153 62 154
rect 62 153 63 154
rect 63 153 64 154
rect 64 153 65 154
rect 215 153 216 154
rect 216 153 217 154
rect 217 153 218 154
rect 218 153 219 154
rect 219 153 220 154
rect 220 153 221 154
rect 221 153 222 154
rect 222 153 223 154
rect 223 153 224 154
rect 224 153 225 154
rect 225 153 226 154
rect 226 153 227 154
rect 15 152 16 153
rect 16 152 17 153
rect 17 152 18 153
rect 18 152 19 153
rect 19 152 20 153
rect 20 152 21 153
rect 21 152 22 153
rect 22 152 23 153
rect 23 152 24 153
rect 24 152 25 153
rect 25 152 26 153
rect 56 152 57 153
rect 57 152 58 153
rect 58 152 59 153
rect 59 152 60 153
rect 60 152 61 153
rect 61 152 62 153
rect 62 152 63 153
rect 63 152 64 153
rect 64 152 65 153
rect 216 152 217 153
rect 217 152 218 153
rect 218 152 219 153
rect 219 152 220 153
rect 220 152 221 153
rect 221 152 222 153
rect 222 152 223 153
rect 223 152 224 153
rect 224 152 225 153
rect 225 152 226 153
rect 226 152 227 153
rect 13 151 14 152
rect 14 151 15 152
rect 15 151 16 152
rect 16 151 17 152
rect 17 151 18 152
rect 18 151 19 152
rect 19 151 20 152
rect 20 151 21 152
rect 21 151 22 152
rect 22 151 23 152
rect 55 151 56 152
rect 56 151 57 152
rect 57 151 58 152
rect 58 151 59 152
rect 59 151 60 152
rect 60 151 61 152
rect 61 151 62 152
rect 62 151 63 152
rect 63 151 64 152
rect 216 151 217 152
rect 217 151 218 152
rect 218 151 219 152
rect 219 151 220 152
rect 220 151 221 152
rect 221 151 222 152
rect 222 151 223 152
rect 223 151 224 152
rect 224 151 225 152
rect 225 151 226 152
rect 226 151 227 152
rect 227 151 228 152
rect 11 150 12 151
rect 12 150 13 151
rect 13 150 14 151
rect 14 150 15 151
rect 15 150 16 151
rect 16 150 17 151
rect 17 150 18 151
rect 18 150 19 151
rect 19 150 20 151
rect 54 150 55 151
rect 55 150 56 151
rect 56 150 57 151
rect 57 150 58 151
rect 58 150 59 151
rect 59 150 60 151
rect 60 150 61 151
rect 61 150 62 151
rect 62 150 63 151
rect 217 150 218 151
rect 218 150 219 151
rect 219 150 220 151
rect 220 150 221 151
rect 221 150 222 151
rect 222 150 223 151
rect 223 150 224 151
rect 224 150 225 151
rect 225 150 226 151
rect 226 150 227 151
rect 227 150 228 151
rect 10 149 11 150
rect 11 149 12 150
rect 12 149 13 150
rect 13 149 14 150
rect 14 149 15 150
rect 15 149 16 150
rect 16 149 17 150
rect 17 149 18 150
rect 18 149 19 150
rect 54 149 55 150
rect 55 149 56 150
rect 56 149 57 150
rect 57 149 58 150
rect 58 149 59 150
rect 59 149 60 150
rect 60 149 61 150
rect 61 149 62 150
rect 62 149 63 150
rect 217 149 218 150
rect 218 149 219 150
rect 219 149 220 150
rect 220 149 221 150
rect 221 149 222 150
rect 222 149 223 150
rect 223 149 224 150
rect 224 149 225 150
rect 225 149 226 150
rect 226 149 227 150
rect 227 149 228 150
rect 9 148 10 149
rect 10 148 11 149
rect 11 148 12 149
rect 12 148 13 149
rect 13 148 14 149
rect 14 148 15 149
rect 52 148 53 149
rect 53 148 54 149
rect 54 148 55 149
rect 55 148 56 149
rect 56 148 57 149
rect 57 148 58 149
rect 58 148 59 149
rect 59 148 60 149
rect 60 148 61 149
rect 61 148 62 149
rect 217 148 218 149
rect 218 148 219 149
rect 219 148 220 149
rect 220 148 221 149
rect 221 148 222 149
rect 222 148 223 149
rect 223 148 224 149
rect 224 148 225 149
rect 225 148 226 149
rect 226 148 227 149
rect 227 148 228 149
rect 228 148 229 149
rect 9 147 10 148
rect 10 147 11 148
rect 11 147 12 148
rect 12 147 13 148
rect 13 147 14 148
rect 51 147 52 148
rect 52 147 53 148
rect 53 147 54 148
rect 54 147 55 148
rect 55 147 56 148
rect 56 147 57 148
rect 57 147 58 148
rect 58 147 59 148
rect 59 147 60 148
rect 219 147 220 148
rect 220 147 221 148
rect 221 147 222 148
rect 222 147 223 148
rect 223 147 224 148
rect 224 147 225 148
rect 225 147 226 148
rect 226 147 227 148
rect 227 147 228 148
rect 228 147 229 148
rect 9 146 10 147
rect 10 146 11 147
rect 11 146 12 147
rect 12 146 13 147
rect 13 146 14 147
rect 14 146 15 147
rect 50 146 51 147
rect 51 146 52 147
rect 52 146 53 147
rect 53 146 54 147
rect 54 146 55 147
rect 55 146 56 147
rect 56 146 57 147
rect 57 146 58 147
rect 58 146 59 147
rect 219 146 220 147
rect 220 146 221 147
rect 221 146 222 147
rect 222 146 223 147
rect 223 146 224 147
rect 224 146 225 147
rect 225 146 226 147
rect 226 146 227 147
rect 227 146 228 147
rect 228 146 229 147
rect 9 145 10 146
rect 10 145 11 146
rect 11 145 12 146
rect 12 145 13 146
rect 13 145 14 146
rect 14 145 15 146
rect 50 145 51 146
rect 51 145 52 146
rect 52 145 53 146
rect 53 145 54 146
rect 54 145 55 146
rect 55 145 56 146
rect 56 145 57 146
rect 57 145 58 146
rect 58 145 59 146
rect 220 145 221 146
rect 221 145 222 146
rect 222 145 223 146
rect 223 145 224 146
rect 224 145 225 146
rect 225 145 226 146
rect 226 145 227 146
rect 227 145 228 146
rect 228 145 229 146
rect 229 145 230 146
rect 9 144 10 145
rect 10 144 11 145
rect 11 144 12 145
rect 12 144 13 145
rect 13 144 14 145
rect 14 144 15 145
rect 50 144 51 145
rect 51 144 52 145
rect 52 144 53 145
rect 53 144 54 145
rect 54 144 55 145
rect 55 144 56 145
rect 56 144 57 145
rect 57 144 58 145
rect 221 144 222 145
rect 222 144 223 145
rect 223 144 224 145
rect 224 144 225 145
rect 225 144 226 145
rect 226 144 227 145
rect 227 144 228 145
rect 228 144 229 145
rect 229 144 230 145
rect 9 143 10 144
rect 10 143 11 144
rect 11 143 12 144
rect 12 143 13 144
rect 13 143 14 144
rect 14 143 15 144
rect 50 143 51 144
rect 51 143 52 144
rect 52 143 53 144
rect 53 143 54 144
rect 54 143 55 144
rect 55 143 56 144
rect 56 143 57 144
rect 221 143 222 144
rect 222 143 223 144
rect 223 143 224 144
rect 224 143 225 144
rect 225 143 226 144
rect 226 143 227 144
rect 227 143 228 144
rect 228 143 229 144
rect 229 143 230 144
rect 9 142 10 143
rect 10 142 11 143
rect 11 142 12 143
rect 12 142 13 143
rect 13 142 14 143
rect 14 142 15 143
rect 15 142 16 143
rect 49 142 50 143
rect 50 142 51 143
rect 51 142 52 143
rect 52 142 53 143
rect 53 142 54 143
rect 54 142 55 143
rect 55 142 56 143
rect 221 142 222 143
rect 222 142 223 143
rect 223 142 224 143
rect 224 142 225 143
rect 225 142 226 143
rect 226 142 227 143
rect 227 142 228 143
rect 228 142 229 143
rect 229 142 230 143
rect 9 141 10 142
rect 10 141 11 142
rect 11 141 12 142
rect 12 141 13 142
rect 13 141 14 142
rect 14 141 15 142
rect 15 141 16 142
rect 16 141 17 142
rect 48 141 49 142
rect 49 141 50 142
rect 50 141 51 142
rect 51 141 52 142
rect 52 141 53 142
rect 53 141 54 142
rect 54 141 55 142
rect 221 141 222 142
rect 222 141 223 142
rect 223 141 224 142
rect 224 141 225 142
rect 225 141 226 142
rect 226 141 227 142
rect 227 141 228 142
rect 228 141 229 142
rect 229 141 230 142
rect 9 140 10 141
rect 10 140 11 141
rect 11 140 12 141
rect 12 140 13 141
rect 13 140 14 141
rect 14 140 15 141
rect 15 140 16 141
rect 16 140 17 141
rect 17 140 18 141
rect 48 140 49 141
rect 49 140 50 141
rect 50 140 51 141
rect 51 140 52 141
rect 52 140 53 141
rect 53 140 54 141
rect 54 140 55 141
rect 223 140 224 141
rect 224 140 225 141
rect 225 140 226 141
rect 226 140 227 141
rect 227 140 228 141
rect 228 140 229 141
rect 229 140 230 141
rect 10 139 11 140
rect 11 139 12 140
rect 12 139 13 140
rect 13 139 14 140
rect 14 139 15 140
rect 15 139 16 140
rect 16 139 17 140
rect 17 139 18 140
rect 47 139 48 140
rect 48 139 49 140
rect 49 139 50 140
rect 50 139 51 140
rect 51 139 52 140
rect 52 139 53 140
rect 53 139 54 140
rect 223 139 224 140
rect 224 139 225 140
rect 225 139 226 140
rect 226 139 227 140
rect 227 139 228 140
rect 228 139 229 140
rect 229 139 230 140
rect 10 138 11 139
rect 11 138 12 139
rect 12 138 13 139
rect 13 138 14 139
rect 14 138 15 139
rect 15 138 16 139
rect 16 138 17 139
rect 17 138 18 139
rect 18 138 19 139
rect 47 138 48 139
rect 48 138 49 139
rect 49 138 50 139
rect 50 138 51 139
rect 51 138 52 139
rect 52 138 53 139
rect 223 138 224 139
rect 224 138 225 139
rect 225 138 226 139
rect 226 138 227 139
rect 227 138 228 139
rect 228 138 229 139
rect 229 138 230 139
rect 10 137 11 138
rect 11 137 12 138
rect 12 137 13 138
rect 13 137 14 138
rect 14 137 15 138
rect 15 137 16 138
rect 16 137 17 138
rect 17 137 18 138
rect 18 137 19 138
rect 47 137 48 138
rect 48 137 49 138
rect 49 137 50 138
rect 50 137 51 138
rect 51 137 52 138
rect 224 137 225 138
rect 225 137 226 138
rect 226 137 227 138
rect 227 137 228 138
rect 228 137 229 138
rect 229 137 230 138
rect 10 136 11 137
rect 11 136 12 137
rect 12 136 13 137
rect 13 136 14 137
rect 14 136 15 137
rect 15 136 16 137
rect 16 136 17 137
rect 17 136 18 137
rect 18 136 19 137
rect 19 136 20 137
rect 46 136 47 137
rect 47 136 48 137
rect 48 136 49 137
rect 49 136 50 137
rect 50 136 51 137
rect 225 136 226 137
rect 226 136 227 137
rect 227 136 228 137
rect 228 136 229 137
rect 229 136 230 137
rect 10 135 11 136
rect 11 135 12 136
rect 12 135 13 136
rect 13 135 14 136
rect 14 135 15 136
rect 15 135 16 136
rect 16 135 17 136
rect 17 135 18 136
rect 18 135 19 136
rect 19 135 20 136
rect 46 135 47 136
rect 47 135 48 136
rect 48 135 49 136
rect 49 135 50 136
rect 50 135 51 136
rect 225 135 226 136
rect 226 135 227 136
rect 227 135 228 136
rect 228 135 229 136
rect 229 135 230 136
rect 11 134 12 135
rect 12 134 13 135
rect 13 134 14 135
rect 14 134 15 135
rect 15 134 16 135
rect 16 134 17 135
rect 17 134 18 135
rect 18 134 19 135
rect 19 134 20 135
rect 20 134 21 135
rect 21 134 22 135
rect 46 134 47 135
rect 47 134 48 135
rect 48 134 49 135
rect 49 134 50 135
rect 50 134 51 135
rect 225 134 226 135
rect 226 134 227 135
rect 227 134 228 135
rect 228 134 229 135
rect 229 134 230 135
rect 230 134 231 135
rect 12 133 13 134
rect 13 133 14 134
rect 14 133 15 134
rect 15 133 16 134
rect 16 133 17 134
rect 17 133 18 134
rect 18 133 19 134
rect 19 133 20 134
rect 20 133 21 134
rect 21 133 22 134
rect 22 133 23 134
rect 45 133 46 134
rect 46 133 47 134
rect 47 133 48 134
rect 48 133 49 134
rect 49 133 50 134
rect 225 133 226 134
rect 226 133 227 134
rect 227 133 228 134
rect 228 133 229 134
rect 229 133 230 134
rect 230 133 231 134
rect 14 132 15 133
rect 15 132 16 133
rect 16 132 17 133
rect 17 132 18 133
rect 18 132 19 133
rect 19 132 20 133
rect 20 132 21 133
rect 21 132 22 133
rect 22 132 23 133
rect 23 132 24 133
rect 45 132 46 133
rect 46 132 47 133
rect 47 132 48 133
rect 48 132 49 133
rect 225 132 226 133
rect 226 132 227 133
rect 227 132 228 133
rect 228 132 229 133
rect 229 132 230 133
rect 230 132 231 133
rect 14 131 15 132
rect 15 131 16 132
rect 16 131 17 132
rect 17 131 18 132
rect 18 131 19 132
rect 19 131 20 132
rect 20 131 21 132
rect 21 131 22 132
rect 22 131 23 132
rect 23 131 24 132
rect 24 131 25 132
rect 44 131 45 132
rect 45 131 46 132
rect 46 131 47 132
rect 47 131 48 132
rect 225 131 226 132
rect 226 131 227 132
rect 227 131 228 132
rect 228 131 229 132
rect 229 131 230 132
rect 230 131 231 132
rect 14 130 15 131
rect 15 130 16 131
rect 16 130 17 131
rect 17 130 18 131
rect 18 130 19 131
rect 19 130 20 131
rect 20 130 21 131
rect 21 130 22 131
rect 22 130 23 131
rect 23 130 24 131
rect 24 130 25 131
rect 25 130 26 131
rect 44 130 45 131
rect 45 130 46 131
rect 46 130 47 131
rect 47 130 48 131
rect 225 130 226 131
rect 226 130 227 131
rect 227 130 228 131
rect 228 130 229 131
rect 229 130 230 131
rect 230 130 231 131
rect 16 129 17 130
rect 17 129 18 130
rect 18 129 19 130
rect 19 129 20 130
rect 20 129 21 130
rect 21 129 22 130
rect 22 129 23 130
rect 23 129 24 130
rect 24 129 25 130
rect 25 129 26 130
rect 26 129 27 130
rect 43 129 44 130
rect 44 129 45 130
rect 45 129 46 130
rect 46 129 47 130
rect 50 129 51 130
rect 51 129 52 130
rect 52 129 53 130
rect 53 129 54 130
rect 54 129 55 130
rect 55 129 56 130
rect 56 129 57 130
rect 57 129 58 130
rect 58 129 59 130
rect 59 129 60 130
rect 60 129 61 130
rect 61 129 62 130
rect 62 129 63 130
rect 64 129 65 130
rect 65 129 66 130
rect 66 129 67 130
rect 67 129 68 130
rect 68 129 69 130
rect 69 129 70 130
rect 70 129 71 130
rect 71 129 72 130
rect 72 129 73 130
rect 73 129 74 130
rect 74 129 75 130
rect 75 129 76 130
rect 226 129 227 130
rect 227 129 228 130
rect 228 129 229 130
rect 229 129 230 130
rect 230 129 231 130
rect 18 128 19 129
rect 19 128 20 129
rect 20 128 21 129
rect 21 128 22 129
rect 22 128 23 129
rect 23 128 24 129
rect 24 128 25 129
rect 25 128 26 129
rect 26 128 27 129
rect 27 128 28 129
rect 42 128 43 129
rect 43 128 44 129
rect 44 128 45 129
rect 45 128 46 129
rect 46 128 47 129
rect 50 128 51 129
rect 51 128 52 129
rect 52 128 53 129
rect 53 128 54 129
rect 54 128 55 129
rect 55 128 56 129
rect 56 128 57 129
rect 57 128 58 129
rect 58 128 59 129
rect 59 128 60 129
rect 60 128 61 129
rect 61 128 62 129
rect 62 128 63 129
rect 64 128 65 129
rect 65 128 66 129
rect 66 128 67 129
rect 67 128 68 129
rect 68 128 69 129
rect 69 128 70 129
rect 70 128 71 129
rect 71 128 72 129
rect 72 128 73 129
rect 73 128 74 129
rect 74 128 75 129
rect 75 128 76 129
rect 226 128 227 129
rect 227 128 228 129
rect 228 128 229 129
rect 229 128 230 129
rect 230 128 231 129
rect 19 127 20 128
rect 20 127 21 128
rect 21 127 22 128
rect 22 127 23 128
rect 23 127 24 128
rect 24 127 25 128
rect 25 127 26 128
rect 26 127 27 128
rect 27 127 28 128
rect 28 127 29 128
rect 29 127 30 128
rect 30 127 31 128
rect 31 127 32 128
rect 41 127 42 128
rect 42 127 43 128
rect 43 127 44 128
rect 44 127 45 128
rect 45 127 46 128
rect 46 127 47 128
rect 52 127 53 128
rect 53 127 54 128
rect 54 127 55 128
rect 55 127 56 128
rect 56 127 57 128
rect 57 127 58 128
rect 58 127 59 128
rect 59 127 60 128
rect 60 127 61 128
rect 67 127 68 128
rect 68 127 69 128
rect 69 127 70 128
rect 70 127 71 128
rect 71 127 72 128
rect 72 127 73 128
rect 73 127 74 128
rect 226 127 227 128
rect 227 127 228 128
rect 228 127 229 128
rect 229 127 230 128
rect 230 127 231 128
rect 22 126 23 127
rect 23 126 24 127
rect 24 126 25 127
rect 25 126 26 127
rect 26 126 27 127
rect 27 126 28 127
rect 28 126 29 127
rect 29 126 30 127
rect 30 126 31 127
rect 31 126 32 127
rect 32 126 33 127
rect 33 126 34 127
rect 34 126 35 127
rect 35 126 36 127
rect 39 126 40 127
rect 40 126 41 127
rect 41 126 42 127
rect 42 126 43 127
rect 43 126 44 127
rect 44 126 45 127
rect 45 126 46 127
rect 54 126 55 127
rect 55 126 56 127
rect 56 126 57 127
rect 57 126 58 127
rect 58 126 59 127
rect 67 126 68 127
rect 68 126 69 127
rect 69 126 70 127
rect 70 126 71 127
rect 71 126 72 127
rect 226 126 227 127
rect 227 126 228 127
rect 228 126 229 127
rect 229 126 230 127
rect 230 126 231 127
rect 24 125 25 126
rect 25 125 26 126
rect 26 125 27 126
rect 27 125 28 126
rect 28 125 29 126
rect 29 125 30 126
rect 30 125 31 126
rect 31 125 32 126
rect 32 125 33 126
rect 33 125 34 126
rect 34 125 35 126
rect 35 125 36 126
rect 36 125 37 126
rect 37 125 38 126
rect 38 125 39 126
rect 39 125 40 126
rect 40 125 41 126
rect 41 125 42 126
rect 42 125 43 126
rect 43 125 44 126
rect 44 125 45 126
rect 54 125 55 126
rect 55 125 56 126
rect 56 125 57 126
rect 57 125 58 126
rect 58 125 59 126
rect 67 125 68 126
rect 68 125 69 126
rect 69 125 70 126
rect 70 125 71 126
rect 227 125 228 126
rect 228 125 229 126
rect 229 125 230 126
rect 230 125 231 126
rect 26 124 27 125
rect 27 124 28 125
rect 28 124 29 125
rect 29 124 30 125
rect 30 124 31 125
rect 31 124 32 125
rect 32 124 33 125
rect 33 124 34 125
rect 34 124 35 125
rect 35 124 36 125
rect 36 124 37 125
rect 37 124 38 125
rect 38 124 39 125
rect 39 124 40 125
rect 40 124 41 125
rect 41 124 42 125
rect 42 124 43 125
rect 43 124 44 125
rect 44 124 45 125
rect 54 124 55 125
rect 55 124 56 125
rect 56 124 57 125
rect 57 124 58 125
rect 58 124 59 125
rect 66 124 67 125
rect 67 124 68 125
rect 68 124 69 125
rect 69 124 70 125
rect 227 124 228 125
rect 228 124 229 125
rect 229 124 230 125
rect 230 124 231 125
rect 28 123 29 124
rect 29 123 30 124
rect 30 123 31 124
rect 31 123 32 124
rect 32 123 33 124
rect 33 123 34 124
rect 34 123 35 124
rect 35 123 36 124
rect 36 123 37 124
rect 37 123 38 124
rect 38 123 39 124
rect 39 123 40 124
rect 40 123 41 124
rect 41 123 42 124
rect 42 123 43 124
rect 43 123 44 124
rect 44 123 45 124
rect 54 123 55 124
rect 55 123 56 124
rect 56 123 57 124
rect 57 123 58 124
rect 58 123 59 124
rect 65 123 66 124
rect 66 123 67 124
rect 67 123 68 124
rect 68 123 69 124
rect 227 123 228 124
rect 228 123 229 124
rect 229 123 230 124
rect 230 123 231 124
rect 30 122 31 123
rect 31 122 32 123
rect 32 122 33 123
rect 33 122 34 123
rect 34 122 35 123
rect 35 122 36 123
rect 36 122 37 123
rect 37 122 38 123
rect 38 122 39 123
rect 39 122 40 123
rect 40 122 41 123
rect 41 122 42 123
rect 42 122 43 123
rect 43 122 44 123
rect 54 122 55 123
rect 55 122 56 123
rect 56 122 57 123
rect 57 122 58 123
rect 58 122 59 123
rect 63 122 64 123
rect 64 122 65 123
rect 65 122 66 123
rect 66 122 67 123
rect 67 122 68 123
rect 227 122 228 123
rect 228 122 229 123
rect 229 122 230 123
rect 230 122 231 123
rect 31 121 32 122
rect 32 121 33 122
rect 33 121 34 122
rect 34 121 35 122
rect 35 121 36 122
rect 36 121 37 122
rect 37 121 38 122
rect 38 121 39 122
rect 39 121 40 122
rect 40 121 41 122
rect 41 121 42 122
rect 42 121 43 122
rect 43 121 44 122
rect 54 121 55 122
rect 55 121 56 122
rect 56 121 57 122
rect 57 121 58 122
rect 58 121 59 122
rect 63 121 64 122
rect 64 121 65 122
rect 65 121 66 122
rect 66 121 67 122
rect 67 121 68 122
rect 227 121 228 122
rect 228 121 229 122
rect 229 121 230 122
rect 230 121 231 122
rect 33 120 34 121
rect 34 120 35 121
rect 35 120 36 121
rect 36 120 37 121
rect 37 120 38 121
rect 38 120 39 121
rect 39 120 40 121
rect 40 120 41 121
rect 41 120 42 121
rect 42 120 43 121
rect 54 120 55 121
rect 55 120 56 121
rect 56 120 57 121
rect 57 120 58 121
rect 58 120 59 121
rect 61 120 62 121
rect 62 120 63 121
rect 63 120 64 121
rect 64 120 65 121
rect 65 120 66 121
rect 66 120 67 121
rect 201 120 202 121
rect 202 120 203 121
rect 203 120 204 121
rect 204 120 205 121
rect 205 120 206 121
rect 206 120 207 121
rect 207 120 208 121
rect 208 120 209 121
rect 209 120 210 121
rect 210 120 211 121
rect 211 120 212 121
rect 212 120 213 121
rect 227 120 228 121
rect 228 120 229 121
rect 229 120 230 121
rect 230 120 231 121
rect 35 119 36 120
rect 36 119 37 120
rect 37 119 38 120
rect 38 119 39 120
rect 39 119 40 120
rect 40 119 41 120
rect 41 119 42 120
rect 42 119 43 120
rect 54 119 55 120
rect 55 119 56 120
rect 56 119 57 120
rect 57 119 58 120
rect 58 119 59 120
rect 60 119 61 120
rect 61 119 62 120
rect 62 119 63 120
rect 63 119 64 120
rect 64 119 65 120
rect 201 119 202 120
rect 202 119 203 120
rect 203 119 204 120
rect 204 119 205 120
rect 205 119 206 120
rect 206 119 207 120
rect 207 119 208 120
rect 208 119 209 120
rect 209 119 210 120
rect 210 119 211 120
rect 211 119 212 120
rect 212 119 213 120
rect 227 119 228 120
rect 228 119 229 120
rect 229 119 230 120
rect 230 119 231 120
rect 37 118 38 119
rect 38 118 39 119
rect 39 118 40 119
rect 40 118 41 119
rect 41 118 42 119
rect 42 118 43 119
rect 54 118 55 119
rect 55 118 56 119
rect 56 118 57 119
rect 57 118 58 119
rect 58 118 59 119
rect 59 118 60 119
rect 60 118 61 119
rect 61 118 62 119
rect 62 118 63 119
rect 63 118 64 119
rect 203 118 204 119
rect 204 118 205 119
rect 205 118 206 119
rect 206 118 207 119
rect 207 118 208 119
rect 208 118 209 119
rect 209 118 210 119
rect 227 118 228 119
rect 228 118 229 119
rect 229 118 230 119
rect 230 118 231 119
rect 38 117 39 118
rect 39 117 40 118
rect 40 117 41 118
rect 41 117 42 118
rect 42 117 43 118
rect 54 117 55 118
rect 55 117 56 118
rect 56 117 57 118
rect 57 117 58 118
rect 58 117 59 118
rect 59 117 60 118
rect 60 117 61 118
rect 61 117 62 118
rect 62 117 63 118
rect 63 117 64 118
rect 204 117 205 118
rect 205 117 206 118
rect 206 117 207 118
rect 207 117 208 118
rect 208 117 209 118
rect 209 117 210 118
rect 227 117 228 118
rect 228 117 229 118
rect 229 117 230 118
rect 230 117 231 118
rect 38 116 39 117
rect 39 116 40 117
rect 40 116 41 117
rect 41 116 42 117
rect 42 116 43 117
rect 54 116 55 117
rect 55 116 56 117
rect 56 116 57 117
rect 57 116 58 117
rect 58 116 59 117
rect 59 116 60 117
rect 60 116 61 117
rect 61 116 62 117
rect 62 116 63 117
rect 63 116 64 117
rect 204 116 205 117
rect 205 116 206 117
rect 206 116 207 117
rect 207 116 208 117
rect 208 116 209 117
rect 209 116 210 117
rect 227 116 228 117
rect 228 116 229 117
rect 229 116 230 117
rect 230 116 231 117
rect 38 115 39 116
rect 39 115 40 116
rect 40 115 41 116
rect 41 115 42 116
rect 42 115 43 116
rect 54 115 55 116
rect 55 115 56 116
rect 56 115 57 116
rect 57 115 58 116
rect 58 115 59 116
rect 59 115 60 116
rect 60 115 61 116
rect 61 115 62 116
rect 62 115 63 116
rect 63 115 64 116
rect 64 115 65 116
rect 204 115 205 116
rect 205 115 206 116
rect 206 115 207 116
rect 207 115 208 116
rect 208 115 209 116
rect 209 115 210 116
rect 227 115 228 116
rect 228 115 229 116
rect 229 115 230 116
rect 230 115 231 116
rect 39 114 40 115
rect 40 114 41 115
rect 41 114 42 115
rect 42 114 43 115
rect 54 114 55 115
rect 55 114 56 115
rect 56 114 57 115
rect 57 114 58 115
rect 58 114 59 115
rect 59 114 60 115
rect 60 114 61 115
rect 61 114 62 115
rect 62 114 63 115
rect 63 114 64 115
rect 64 114 65 115
rect 65 114 66 115
rect 66 114 67 115
rect 204 114 205 115
rect 205 114 206 115
rect 206 114 207 115
rect 207 114 208 115
rect 208 114 209 115
rect 209 114 210 115
rect 227 114 228 115
rect 228 114 229 115
rect 229 114 230 115
rect 230 114 231 115
rect 40 113 41 114
rect 41 113 42 114
rect 54 113 55 114
rect 55 113 56 114
rect 56 113 57 114
rect 57 113 58 114
rect 58 113 59 114
rect 60 113 61 114
rect 61 113 62 114
rect 62 113 63 114
rect 63 113 64 114
rect 64 113 65 114
rect 65 113 66 114
rect 66 113 67 114
rect 67 113 68 114
rect 204 113 205 114
rect 205 113 206 114
rect 206 113 207 114
rect 207 113 208 114
rect 208 113 209 114
rect 209 113 210 114
rect 227 113 228 114
rect 228 113 229 114
rect 229 113 230 114
rect 230 113 231 114
rect 40 112 41 113
rect 41 112 42 113
rect 54 112 55 113
rect 55 112 56 113
rect 56 112 57 113
rect 57 112 58 113
rect 58 112 59 113
rect 61 112 62 113
rect 62 112 63 113
rect 63 112 64 113
rect 64 112 65 113
rect 65 112 66 113
rect 66 112 67 113
rect 67 112 68 113
rect 82 112 83 113
rect 83 112 84 113
rect 204 112 205 113
rect 205 112 206 113
rect 206 112 207 113
rect 207 112 208 113
rect 208 112 209 113
rect 209 112 210 113
rect 227 112 228 113
rect 228 112 229 113
rect 229 112 230 113
rect 230 112 231 113
rect 40 111 41 112
rect 41 111 42 112
rect 54 111 55 112
rect 55 111 56 112
rect 56 111 57 112
rect 57 111 58 112
rect 58 111 59 112
rect 62 111 63 112
rect 63 111 64 112
rect 64 111 65 112
rect 65 111 66 112
rect 66 111 67 112
rect 67 111 68 112
rect 68 111 69 112
rect 82 111 83 112
rect 83 111 84 112
rect 84 111 85 112
rect 204 111 205 112
rect 205 111 206 112
rect 206 111 207 112
rect 207 111 208 112
rect 208 111 209 112
rect 209 111 210 112
rect 227 111 228 112
rect 228 111 229 112
rect 229 111 230 112
rect 230 111 231 112
rect 54 110 55 111
rect 55 110 56 111
rect 56 110 57 111
rect 57 110 58 111
rect 58 110 59 111
rect 63 110 64 111
rect 64 110 65 111
rect 65 110 66 111
rect 66 110 67 111
rect 67 110 68 111
rect 68 110 69 111
rect 81 110 82 111
rect 82 110 83 111
rect 83 110 84 111
rect 84 110 85 111
rect 204 110 205 111
rect 205 110 206 111
rect 206 110 207 111
rect 207 110 208 111
rect 208 110 209 111
rect 209 110 210 111
rect 227 110 228 111
rect 228 110 229 111
rect 229 110 230 111
rect 230 110 231 111
rect 40 109 41 110
rect 41 109 42 110
rect 54 109 55 110
rect 55 109 56 110
rect 56 109 57 110
rect 57 109 58 110
rect 58 109 59 110
rect 63 109 64 110
rect 64 109 65 110
rect 65 109 66 110
rect 66 109 67 110
rect 67 109 68 110
rect 68 109 69 110
rect 69 109 70 110
rect 70 109 71 110
rect 81 109 82 110
rect 82 109 83 110
rect 83 109 84 110
rect 84 109 85 110
rect 204 109 205 110
rect 205 109 206 110
rect 206 109 207 110
rect 207 109 208 110
rect 208 109 209 110
rect 209 109 210 110
rect 227 109 228 110
rect 228 109 229 110
rect 229 109 230 110
rect 230 109 231 110
rect 40 108 41 109
rect 41 108 42 109
rect 54 108 55 109
rect 55 108 56 109
rect 56 108 57 109
rect 57 108 58 109
rect 58 108 59 109
rect 64 108 65 109
rect 65 108 66 109
rect 66 108 67 109
rect 67 108 68 109
rect 68 108 69 109
rect 69 108 70 109
rect 70 108 71 109
rect 71 108 72 109
rect 80 108 81 109
rect 81 108 82 109
rect 82 108 83 109
rect 83 108 84 109
rect 84 108 85 109
rect 85 108 86 109
rect 204 108 205 109
rect 205 108 206 109
rect 206 108 207 109
rect 207 108 208 109
rect 208 108 209 109
rect 209 108 210 109
rect 227 108 228 109
rect 228 108 229 109
rect 229 108 230 109
rect 230 108 231 109
rect 40 107 41 108
rect 41 107 42 108
rect 54 107 55 108
rect 55 107 56 108
rect 56 107 57 108
rect 57 107 58 108
rect 58 107 59 108
rect 65 107 66 108
rect 66 107 67 108
rect 67 107 68 108
rect 68 107 69 108
rect 69 107 70 108
rect 70 107 71 108
rect 71 107 72 108
rect 80 107 81 108
rect 81 107 82 108
rect 82 107 83 108
rect 83 107 84 108
rect 84 107 85 108
rect 85 107 86 108
rect 86 107 87 108
rect 204 107 205 108
rect 205 107 206 108
rect 206 107 207 108
rect 207 107 208 108
rect 208 107 209 108
rect 209 107 210 108
rect 227 107 228 108
rect 228 107 229 108
rect 229 107 230 108
rect 230 107 231 108
rect 40 106 41 107
rect 41 106 42 107
rect 54 106 55 107
rect 55 106 56 107
rect 56 106 57 107
rect 57 106 58 107
rect 58 106 59 107
rect 66 106 67 107
rect 67 106 68 107
rect 68 106 69 107
rect 69 106 70 107
rect 70 106 71 107
rect 71 106 72 107
rect 72 106 73 107
rect 79 106 80 107
rect 80 106 81 107
rect 81 106 82 107
rect 82 106 83 107
rect 83 106 84 107
rect 84 106 85 107
rect 85 106 86 107
rect 86 106 87 107
rect 204 106 205 107
rect 205 106 206 107
rect 206 106 207 107
rect 207 106 208 107
rect 208 106 209 107
rect 209 106 210 107
rect 227 106 228 107
rect 228 106 229 107
rect 229 106 230 107
rect 230 106 231 107
rect 40 105 41 106
rect 41 105 42 106
rect 54 105 55 106
rect 55 105 56 106
rect 56 105 57 106
rect 57 105 58 106
rect 58 105 59 106
rect 67 105 68 106
rect 68 105 69 106
rect 69 105 70 106
rect 70 105 71 106
rect 71 105 72 106
rect 72 105 73 106
rect 73 105 74 106
rect 79 105 80 106
rect 80 105 81 106
rect 81 105 82 106
rect 82 105 83 106
rect 83 105 84 106
rect 84 105 85 106
rect 85 105 86 106
rect 86 105 87 106
rect 87 105 88 106
rect 204 105 205 106
rect 205 105 206 106
rect 206 105 207 106
rect 207 105 208 106
rect 208 105 209 106
rect 209 105 210 106
rect 226 105 227 106
rect 227 105 228 106
rect 228 105 229 106
rect 229 105 230 106
rect 40 104 41 105
rect 41 104 42 105
rect 54 104 55 105
rect 55 104 56 105
rect 56 104 57 105
rect 57 104 58 105
rect 58 104 59 105
rect 67 104 68 105
rect 68 104 69 105
rect 69 104 70 105
rect 70 104 71 105
rect 71 104 72 105
rect 72 104 73 105
rect 73 104 74 105
rect 74 104 75 105
rect 79 104 80 105
rect 80 104 81 105
rect 81 104 82 105
rect 82 104 83 105
rect 83 104 84 105
rect 84 104 85 105
rect 85 104 86 105
rect 86 104 87 105
rect 87 104 88 105
rect 204 104 205 105
rect 205 104 206 105
rect 206 104 207 105
rect 207 104 208 105
rect 208 104 209 105
rect 209 104 210 105
rect 226 104 227 105
rect 227 104 228 105
rect 228 104 229 105
rect 229 104 230 105
rect 40 103 41 104
rect 41 103 42 104
rect 54 103 55 104
rect 55 103 56 104
rect 56 103 57 104
rect 57 103 58 104
rect 58 103 59 104
rect 68 103 69 104
rect 69 103 70 104
rect 70 103 71 104
rect 71 103 72 104
rect 72 103 73 104
rect 73 103 74 104
rect 74 103 75 104
rect 75 103 76 104
rect 79 103 80 104
rect 80 103 81 104
rect 81 103 82 104
rect 83 103 84 104
rect 84 103 85 104
rect 85 103 86 104
rect 86 103 87 104
rect 87 103 88 104
rect 204 103 205 104
rect 205 103 206 104
rect 206 103 207 104
rect 207 103 208 104
rect 208 103 209 104
rect 209 103 210 104
rect 226 103 227 104
rect 227 103 228 104
rect 228 103 229 104
rect 229 103 230 104
rect 39 102 40 103
rect 40 102 41 103
rect 41 102 42 103
rect 50 102 51 103
rect 51 102 52 103
rect 52 102 53 103
rect 53 102 54 103
rect 54 102 55 103
rect 55 102 56 103
rect 56 102 57 103
rect 57 102 58 103
rect 58 102 59 103
rect 59 102 60 103
rect 60 102 61 103
rect 61 102 62 103
rect 66 102 67 103
rect 67 102 68 103
rect 68 102 69 103
rect 69 102 70 103
rect 70 102 71 103
rect 71 102 72 103
rect 72 102 73 103
rect 73 102 74 103
rect 74 102 75 103
rect 75 102 76 103
rect 76 102 77 103
rect 77 102 78 103
rect 78 102 79 103
rect 79 102 80 103
rect 80 102 81 103
rect 81 102 82 103
rect 83 102 84 103
rect 84 102 85 103
rect 85 102 86 103
rect 86 102 87 103
rect 87 102 88 103
rect 204 102 205 103
rect 205 102 206 103
rect 206 102 207 103
rect 207 102 208 103
rect 208 102 209 103
rect 209 102 210 103
rect 226 102 227 103
rect 227 102 228 103
rect 228 102 229 103
rect 229 102 230 103
rect 39 101 40 102
rect 40 101 41 102
rect 41 101 42 102
rect 50 101 51 102
rect 51 101 52 102
rect 52 101 53 102
rect 53 101 54 102
rect 54 101 55 102
rect 55 101 56 102
rect 56 101 57 102
rect 57 101 58 102
rect 58 101 59 102
rect 59 101 60 102
rect 60 101 61 102
rect 61 101 62 102
rect 65 101 66 102
rect 66 101 67 102
rect 67 101 68 102
rect 68 101 69 102
rect 69 101 70 102
rect 70 101 71 102
rect 71 101 72 102
rect 72 101 73 102
rect 73 101 74 102
rect 74 101 75 102
rect 75 101 76 102
rect 76 101 77 102
rect 77 101 78 102
rect 78 101 79 102
rect 79 101 80 102
rect 80 101 81 102
rect 83 101 84 102
rect 84 101 85 102
rect 85 101 86 102
rect 86 101 87 102
rect 87 101 88 102
rect 204 101 205 102
rect 205 101 206 102
rect 206 101 207 102
rect 207 101 208 102
rect 208 101 209 102
rect 209 101 210 102
rect 226 101 227 102
rect 227 101 228 102
rect 228 101 229 102
rect 229 101 230 102
rect 39 100 40 101
rect 40 100 41 101
rect 41 100 42 101
rect 51 100 52 101
rect 52 100 53 101
rect 53 100 54 101
rect 54 100 55 101
rect 55 100 56 101
rect 56 100 57 101
rect 57 100 58 101
rect 58 100 59 101
rect 59 100 60 101
rect 60 100 61 101
rect 65 100 66 101
rect 66 100 67 101
rect 67 100 68 101
rect 68 100 69 101
rect 69 100 70 101
rect 70 100 71 101
rect 71 100 72 101
rect 72 100 73 101
rect 73 100 74 101
rect 74 100 75 101
rect 75 100 76 101
rect 76 100 77 101
rect 77 100 78 101
rect 78 100 79 101
rect 79 100 80 101
rect 80 100 81 101
rect 83 100 84 101
rect 84 100 85 101
rect 85 100 86 101
rect 86 100 87 101
rect 87 100 88 101
rect 88 100 89 101
rect 177 100 178 101
rect 178 100 179 101
rect 179 100 180 101
rect 180 100 181 101
rect 181 100 182 101
rect 182 100 183 101
rect 183 100 184 101
rect 184 100 185 101
rect 185 100 186 101
rect 186 100 187 101
rect 187 100 188 101
rect 188 100 189 101
rect 189 100 190 101
rect 190 100 191 101
rect 191 100 192 101
rect 192 100 193 101
rect 193 100 194 101
rect 194 100 195 101
rect 195 100 196 101
rect 196 100 197 101
rect 197 100 198 101
rect 198 100 199 101
rect 199 100 200 101
rect 200 100 201 101
rect 204 100 205 101
rect 205 100 206 101
rect 206 100 207 101
rect 207 100 208 101
rect 208 100 209 101
rect 209 100 210 101
rect 225 100 226 101
rect 226 100 227 101
rect 227 100 228 101
rect 228 100 229 101
rect 229 100 230 101
rect 38 99 39 100
rect 39 99 40 100
rect 40 99 41 100
rect 41 99 42 100
rect 77 99 78 100
rect 78 99 79 100
rect 79 99 80 100
rect 84 99 85 100
rect 85 99 86 100
rect 86 99 87 100
rect 87 99 88 100
rect 88 99 89 100
rect 89 99 90 100
rect 177 99 178 100
rect 178 99 179 100
rect 179 99 180 100
rect 180 99 181 100
rect 181 99 182 100
rect 182 99 183 100
rect 183 99 184 100
rect 184 99 185 100
rect 185 99 186 100
rect 186 99 187 100
rect 187 99 188 100
rect 188 99 189 100
rect 189 99 190 100
rect 190 99 191 100
rect 191 99 192 100
rect 192 99 193 100
rect 193 99 194 100
rect 194 99 195 100
rect 195 99 196 100
rect 196 99 197 100
rect 197 99 198 100
rect 198 99 199 100
rect 199 99 200 100
rect 200 99 201 100
rect 204 99 205 100
rect 205 99 206 100
rect 206 99 207 100
rect 207 99 208 100
rect 208 99 209 100
rect 209 99 210 100
rect 225 99 226 100
rect 226 99 227 100
rect 227 99 228 100
rect 228 99 229 100
rect 229 99 230 100
rect 38 98 39 99
rect 39 98 40 99
rect 40 98 41 99
rect 41 98 42 99
rect 76 98 77 99
rect 77 98 78 99
rect 78 98 79 99
rect 79 98 80 99
rect 84 98 85 99
rect 85 98 86 99
rect 86 98 87 99
rect 87 98 88 99
rect 88 98 89 99
rect 89 98 90 99
rect 177 98 178 99
rect 178 98 179 99
rect 179 98 180 99
rect 180 98 181 99
rect 181 98 182 99
rect 182 98 183 99
rect 183 98 184 99
rect 184 98 185 99
rect 185 98 186 99
rect 186 98 187 99
rect 187 98 188 99
rect 188 98 189 99
rect 189 98 190 99
rect 190 98 191 99
rect 191 98 192 99
rect 192 98 193 99
rect 193 98 194 99
rect 194 98 195 99
rect 195 98 196 99
rect 196 98 197 99
rect 197 98 198 99
rect 198 98 199 99
rect 199 98 200 99
rect 204 98 205 99
rect 205 98 206 99
rect 206 98 207 99
rect 207 98 208 99
rect 208 98 209 99
rect 209 98 210 99
rect 225 98 226 99
rect 226 98 227 99
rect 227 98 228 99
rect 228 98 229 99
rect 229 98 230 99
rect 38 97 39 98
rect 39 97 40 98
rect 40 97 41 98
rect 41 97 42 98
rect 42 97 43 98
rect 76 97 77 98
rect 77 97 78 98
rect 78 97 79 98
rect 79 97 80 98
rect 85 97 86 98
rect 86 97 87 98
rect 87 97 88 98
rect 88 97 89 98
rect 89 97 90 98
rect 177 97 178 98
rect 178 97 179 98
rect 179 97 180 98
rect 180 97 181 98
rect 181 97 182 98
rect 186 97 187 98
rect 187 97 188 98
rect 188 97 189 98
rect 189 97 190 98
rect 190 97 191 98
rect 196 97 197 98
rect 197 97 198 98
rect 198 97 199 98
rect 199 97 200 98
rect 204 97 205 98
rect 205 97 206 98
rect 206 97 207 98
rect 207 97 208 98
rect 208 97 209 98
rect 209 97 210 98
rect 225 97 226 98
rect 226 97 227 98
rect 227 97 228 98
rect 228 97 229 98
rect 229 97 230 98
rect 38 96 39 97
rect 39 96 40 97
rect 40 96 41 97
rect 41 96 42 97
rect 42 96 43 97
rect 76 96 77 97
rect 77 96 78 97
rect 78 96 79 97
rect 79 96 80 97
rect 85 96 86 97
rect 86 96 87 97
rect 87 96 88 97
rect 88 96 89 97
rect 89 96 90 97
rect 90 96 91 97
rect 176 96 177 97
rect 177 96 178 97
rect 178 96 179 97
rect 179 96 180 97
rect 180 96 181 97
rect 185 96 186 97
rect 186 96 187 97
rect 187 96 188 97
rect 188 96 189 97
rect 189 96 190 97
rect 190 96 191 97
rect 197 96 198 97
rect 198 96 199 97
rect 199 96 200 97
rect 204 96 205 97
rect 205 96 206 97
rect 206 96 207 97
rect 207 96 208 97
rect 208 96 209 97
rect 209 96 210 97
rect 225 96 226 97
rect 226 96 227 97
rect 227 96 228 97
rect 228 96 229 97
rect 229 96 230 97
rect 38 95 39 96
rect 39 95 40 96
rect 40 95 41 96
rect 41 95 42 96
rect 42 95 43 96
rect 75 95 76 96
rect 76 95 77 96
rect 77 95 78 96
rect 78 95 79 96
rect 79 95 80 96
rect 81 95 82 96
rect 82 95 83 96
rect 83 95 84 96
rect 84 95 85 96
rect 85 95 86 96
rect 86 95 87 96
rect 87 95 88 96
rect 88 95 89 96
rect 89 95 90 96
rect 90 95 91 96
rect 176 95 177 96
rect 177 95 178 96
rect 178 95 179 96
rect 179 95 180 96
rect 185 95 186 96
rect 186 95 187 96
rect 187 95 188 96
rect 188 95 189 96
rect 189 95 190 96
rect 190 95 191 96
rect 197 95 198 96
rect 198 95 199 96
rect 199 95 200 96
rect 200 95 201 96
rect 204 95 205 96
rect 205 95 206 96
rect 206 95 207 96
rect 207 95 208 96
rect 208 95 209 96
rect 209 95 210 96
rect 225 95 226 96
rect 226 95 227 96
rect 227 95 228 96
rect 228 95 229 96
rect 229 95 230 96
rect 38 94 39 95
rect 39 94 40 95
rect 40 94 41 95
rect 41 94 42 95
rect 42 94 43 95
rect 75 94 76 95
rect 76 94 77 95
rect 77 94 78 95
rect 78 94 79 95
rect 79 94 80 95
rect 80 94 81 95
rect 81 94 82 95
rect 82 94 83 95
rect 83 94 84 95
rect 84 94 85 95
rect 85 94 86 95
rect 86 94 87 95
rect 87 94 88 95
rect 88 94 89 95
rect 89 94 90 95
rect 90 94 91 95
rect 91 94 92 95
rect 177 94 178 95
rect 178 94 179 95
rect 179 94 180 95
rect 186 94 187 95
rect 187 94 188 95
rect 188 94 189 95
rect 189 94 190 95
rect 190 94 191 95
rect 197 94 198 95
rect 198 94 199 95
rect 199 94 200 95
rect 200 94 201 95
rect 204 94 205 95
rect 205 94 206 95
rect 206 94 207 95
rect 207 94 208 95
rect 208 94 209 95
rect 209 94 210 95
rect 224 94 225 95
rect 225 94 226 95
rect 226 94 227 95
rect 227 94 228 95
rect 228 94 229 95
rect 38 93 39 94
rect 39 93 40 94
rect 40 93 41 94
rect 41 93 42 94
rect 42 93 43 94
rect 75 93 76 94
rect 76 93 77 94
rect 77 93 78 94
rect 78 93 79 94
rect 79 93 80 94
rect 80 93 81 94
rect 81 93 82 94
rect 82 93 83 94
rect 83 93 84 94
rect 84 93 85 94
rect 85 93 86 94
rect 86 93 87 94
rect 87 93 88 94
rect 88 93 89 94
rect 89 93 90 94
rect 90 93 91 94
rect 91 93 92 94
rect 177 93 178 94
rect 178 93 179 94
rect 186 93 187 94
rect 187 93 188 94
rect 188 93 189 94
rect 189 93 190 94
rect 190 93 191 94
rect 197 93 198 94
rect 198 93 199 94
rect 199 93 200 94
rect 201 93 202 94
rect 202 93 203 94
rect 203 93 204 94
rect 204 93 205 94
rect 205 93 206 94
rect 206 93 207 94
rect 207 93 208 94
rect 208 93 209 94
rect 209 93 210 94
rect 210 93 211 94
rect 211 93 212 94
rect 212 93 213 94
rect 224 93 225 94
rect 225 93 226 94
rect 226 93 227 94
rect 227 93 228 94
rect 228 93 229 94
rect 38 92 39 93
rect 39 92 40 93
rect 40 92 41 93
rect 41 92 42 93
rect 42 92 43 93
rect 74 92 75 93
rect 75 92 76 93
rect 76 92 77 93
rect 77 92 78 93
rect 87 92 88 93
rect 88 92 89 93
rect 89 92 90 93
rect 90 92 91 93
rect 91 92 92 93
rect 185 92 186 93
rect 186 92 187 93
rect 187 92 188 93
rect 188 92 189 93
rect 189 92 190 93
rect 190 92 191 93
rect 201 92 202 93
rect 202 92 203 93
rect 203 92 204 93
rect 204 92 205 93
rect 205 92 206 93
rect 206 92 207 93
rect 207 92 208 93
rect 208 92 209 93
rect 209 92 210 93
rect 210 92 211 93
rect 211 92 212 93
rect 212 92 213 93
rect 223 92 224 93
rect 224 92 225 93
rect 225 92 226 93
rect 226 92 227 93
rect 227 92 228 93
rect 228 92 229 93
rect 38 91 39 92
rect 39 91 40 92
rect 40 91 41 92
rect 41 91 42 92
rect 42 91 43 92
rect 74 91 75 92
rect 75 91 76 92
rect 76 91 77 92
rect 87 91 88 92
rect 88 91 89 92
rect 89 91 90 92
rect 90 91 91 92
rect 91 91 92 92
rect 185 91 186 92
rect 186 91 187 92
rect 187 91 188 92
rect 188 91 189 92
rect 189 91 190 92
rect 190 91 191 92
rect 201 91 202 92
rect 203 91 204 92
rect 204 91 205 92
rect 205 91 206 92
rect 206 91 207 92
rect 209 91 210 92
rect 210 91 211 92
rect 211 91 212 92
rect 223 91 224 92
rect 224 91 225 92
rect 225 91 226 92
rect 226 91 227 92
rect 227 91 228 92
rect 228 91 229 92
rect 39 90 40 91
rect 40 90 41 91
rect 41 90 42 91
rect 42 90 43 91
rect 43 90 44 91
rect 74 90 75 91
rect 75 90 76 91
rect 76 90 77 91
rect 87 90 88 91
rect 88 90 89 91
rect 89 90 90 91
rect 90 90 91 91
rect 91 90 92 91
rect 92 90 93 91
rect 186 90 187 91
rect 187 90 188 91
rect 188 90 189 91
rect 189 90 190 91
rect 190 90 191 91
rect 223 90 224 91
rect 224 90 225 91
rect 225 90 226 91
rect 226 90 227 91
rect 227 90 228 91
rect 39 89 40 90
rect 40 89 41 90
rect 41 89 42 90
rect 42 89 43 90
rect 43 89 44 90
rect 73 89 74 90
rect 74 89 75 90
rect 75 89 76 90
rect 76 89 77 90
rect 87 89 88 90
rect 88 89 89 90
rect 89 89 90 90
rect 90 89 91 90
rect 91 89 92 90
rect 92 89 93 90
rect 185 89 186 90
rect 186 89 187 90
rect 187 89 188 90
rect 188 89 189 90
rect 189 89 190 90
rect 190 89 191 90
rect 222 89 223 90
rect 223 89 224 90
rect 224 89 225 90
rect 225 89 226 90
rect 226 89 227 90
rect 227 89 228 90
rect 39 88 40 89
rect 40 88 41 89
rect 41 88 42 89
rect 42 88 43 89
rect 43 88 44 89
rect 73 88 74 89
rect 74 88 75 89
rect 75 88 76 89
rect 88 88 89 89
rect 89 88 90 89
rect 90 88 91 89
rect 91 88 92 89
rect 92 88 93 89
rect 93 88 94 89
rect 96 88 97 89
rect 97 88 98 89
rect 98 88 99 89
rect 185 88 186 89
rect 186 88 187 89
rect 187 88 188 89
rect 188 88 189 89
rect 189 88 190 89
rect 190 88 191 89
rect 222 88 223 89
rect 223 88 224 89
rect 224 88 225 89
rect 225 88 226 89
rect 226 88 227 89
rect 227 88 228 89
rect 39 87 40 88
rect 40 87 41 88
rect 41 87 42 88
rect 42 87 43 88
rect 43 87 44 88
rect 72 87 73 88
rect 73 87 74 88
rect 74 87 75 88
rect 75 87 76 88
rect 88 87 89 88
rect 89 87 90 88
rect 90 87 91 88
rect 91 87 92 88
rect 92 87 93 88
rect 93 87 94 88
rect 96 87 97 88
rect 97 87 98 88
rect 98 87 99 88
rect 186 87 187 88
rect 187 87 188 88
rect 188 87 189 88
rect 189 87 190 88
rect 190 87 191 88
rect 221 87 222 88
rect 222 87 223 88
rect 223 87 224 88
rect 224 87 225 88
rect 225 87 226 88
rect 226 87 227 88
rect 40 86 41 87
rect 41 86 42 87
rect 42 86 43 87
rect 43 86 44 87
rect 44 86 45 87
rect 71 86 72 87
rect 72 86 73 87
rect 73 86 74 87
rect 74 86 75 87
rect 75 86 76 87
rect 88 86 89 87
rect 89 86 90 87
rect 90 86 91 87
rect 91 86 92 87
rect 92 86 93 87
rect 93 86 94 87
rect 94 86 95 87
rect 95 86 96 87
rect 96 86 97 87
rect 97 86 98 87
rect 98 86 99 87
rect 99 86 100 87
rect 185 86 186 87
rect 186 86 187 87
rect 187 86 188 87
rect 188 86 189 87
rect 189 86 190 87
rect 190 86 191 87
rect 221 86 222 87
rect 222 86 223 87
rect 223 86 224 87
rect 224 86 225 87
rect 225 86 226 87
rect 226 86 227 87
rect 40 85 41 86
rect 41 85 42 86
rect 42 85 43 86
rect 43 85 44 86
rect 44 85 45 86
rect 70 85 71 86
rect 71 85 72 86
rect 72 85 73 86
rect 73 85 74 86
rect 74 85 75 86
rect 75 85 76 86
rect 76 85 77 86
rect 77 85 78 86
rect 86 85 87 86
rect 87 85 88 86
rect 88 85 89 86
rect 89 85 90 86
rect 90 85 91 86
rect 91 85 92 86
rect 92 85 93 86
rect 93 85 94 86
rect 94 85 95 86
rect 95 85 96 86
rect 96 85 97 86
rect 97 85 98 86
rect 98 85 99 86
rect 99 85 100 86
rect 154 85 155 86
rect 155 85 156 86
rect 156 85 157 86
rect 157 85 158 86
rect 158 85 159 86
rect 159 85 160 86
rect 160 85 161 86
rect 161 85 162 86
rect 162 85 163 86
rect 163 85 164 86
rect 164 85 165 86
rect 165 85 166 86
rect 166 85 167 86
rect 167 85 168 86
rect 168 85 169 86
rect 169 85 170 86
rect 170 85 171 86
rect 171 85 172 86
rect 172 85 173 86
rect 173 85 174 86
rect 174 85 175 86
rect 186 85 187 86
rect 187 85 188 86
rect 188 85 189 86
rect 189 85 190 86
rect 190 85 191 86
rect 221 85 222 86
rect 222 85 223 86
rect 223 85 224 86
rect 224 85 225 86
rect 225 85 226 86
rect 226 85 227 86
rect 40 84 41 85
rect 41 84 42 85
rect 42 84 43 85
rect 43 84 44 85
rect 44 84 45 85
rect 70 84 71 85
rect 71 84 72 85
rect 72 84 73 85
rect 73 84 74 85
rect 74 84 75 85
rect 75 84 76 85
rect 76 84 77 85
rect 77 84 78 85
rect 86 84 87 85
rect 87 84 88 85
rect 88 84 89 85
rect 89 84 90 85
rect 90 84 91 85
rect 91 84 92 85
rect 92 84 93 85
rect 93 84 94 85
rect 94 84 95 85
rect 95 84 96 85
rect 96 84 97 85
rect 97 84 98 85
rect 98 84 99 85
rect 99 84 100 85
rect 154 84 155 85
rect 155 84 156 85
rect 156 84 157 85
rect 157 84 158 85
rect 158 84 159 85
rect 159 84 160 85
rect 160 84 161 85
rect 161 84 162 85
rect 162 84 163 85
rect 163 84 164 85
rect 164 84 165 85
rect 165 84 166 85
rect 166 84 167 85
rect 167 84 168 85
rect 168 84 169 85
rect 169 84 170 85
rect 170 84 171 85
rect 171 84 172 85
rect 172 84 173 85
rect 173 84 174 85
rect 174 84 175 85
rect 185 84 186 85
rect 186 84 187 85
rect 187 84 188 85
rect 188 84 189 85
rect 189 84 190 85
rect 190 84 191 85
rect 220 84 221 85
rect 221 84 222 85
rect 222 84 223 85
rect 223 84 224 85
rect 224 84 225 85
rect 225 84 226 85
rect 40 83 41 84
rect 41 83 42 84
rect 42 83 43 84
rect 43 83 44 84
rect 44 83 45 84
rect 71 83 72 84
rect 72 83 73 84
rect 73 83 74 84
rect 74 83 75 84
rect 75 83 76 84
rect 76 83 77 84
rect 77 83 78 84
rect 87 83 88 84
rect 88 83 89 84
rect 89 83 90 84
rect 90 83 91 84
rect 91 83 92 84
rect 92 83 93 84
rect 93 83 94 84
rect 94 83 95 84
rect 95 83 96 84
rect 96 83 97 84
rect 97 83 98 84
rect 98 83 99 84
rect 99 83 100 84
rect 154 83 155 84
rect 155 83 156 84
rect 156 83 157 84
rect 157 83 158 84
rect 158 83 159 84
rect 159 83 160 84
rect 160 83 161 84
rect 161 83 162 84
rect 162 83 163 84
rect 163 83 164 84
rect 164 83 165 84
rect 165 83 166 84
rect 166 83 167 84
rect 167 83 168 84
rect 168 83 169 84
rect 169 83 170 84
rect 170 83 171 84
rect 171 83 172 84
rect 172 83 173 84
rect 173 83 174 84
rect 174 83 175 84
rect 185 83 186 84
rect 186 83 187 84
rect 187 83 188 84
rect 188 83 189 84
rect 189 83 190 84
rect 190 83 191 84
rect 220 83 221 84
rect 221 83 222 84
rect 222 83 223 84
rect 223 83 224 84
rect 224 83 225 84
rect 225 83 226 84
rect 41 82 42 83
rect 42 82 43 83
rect 43 82 44 83
rect 44 82 45 83
rect 45 82 46 83
rect 95 82 96 83
rect 96 82 97 83
rect 97 82 98 83
rect 98 82 99 83
rect 99 82 100 83
rect 155 82 156 83
rect 156 82 157 83
rect 157 82 158 83
rect 158 82 159 83
rect 159 82 160 83
rect 160 82 161 83
rect 161 82 162 83
rect 162 82 163 83
rect 163 82 164 83
rect 164 82 165 83
rect 165 82 166 83
rect 166 82 167 83
rect 167 82 168 83
rect 168 82 169 83
rect 169 82 170 83
rect 170 82 171 83
rect 171 82 172 83
rect 172 82 173 83
rect 173 82 174 83
rect 174 82 175 83
rect 186 82 187 83
rect 187 82 188 83
rect 188 82 189 83
rect 189 82 190 83
rect 190 82 191 83
rect 220 82 221 83
rect 221 82 222 83
rect 222 82 223 83
rect 223 82 224 83
rect 224 82 225 83
rect 225 82 226 83
rect 41 81 42 82
rect 42 81 43 82
rect 43 81 44 82
rect 44 81 45 82
rect 45 81 46 82
rect 94 81 95 82
rect 95 81 96 82
rect 96 81 97 82
rect 97 81 98 82
rect 98 81 99 82
rect 99 81 100 82
rect 100 81 101 82
rect 124 81 125 82
rect 125 81 126 82
rect 156 81 157 82
rect 157 81 158 82
rect 158 81 159 82
rect 159 81 160 82
rect 160 81 161 82
rect 161 81 162 82
rect 171 81 172 82
rect 172 81 173 82
rect 173 81 174 82
rect 174 81 175 82
rect 185 81 186 82
rect 186 81 187 82
rect 187 81 188 82
rect 188 81 189 82
rect 189 81 190 82
rect 190 81 191 82
rect 219 81 220 82
rect 220 81 221 82
rect 221 81 222 82
rect 222 81 223 82
rect 223 81 224 82
rect 224 81 225 82
rect 225 81 226 82
rect 41 80 42 81
rect 42 80 43 81
rect 43 80 44 81
rect 44 80 45 81
rect 45 80 46 81
rect 46 80 47 81
rect 94 80 95 81
rect 95 80 96 81
rect 96 80 97 81
rect 97 80 98 81
rect 98 80 99 81
rect 99 80 100 81
rect 100 80 101 81
rect 101 80 102 81
rect 123 80 124 81
rect 124 80 125 81
rect 125 80 126 81
rect 126 80 127 81
rect 156 80 157 81
rect 157 80 158 81
rect 158 80 159 81
rect 159 80 160 81
rect 160 80 161 81
rect 161 80 162 81
rect 162 80 163 81
rect 163 80 164 81
rect 172 80 173 81
rect 173 80 174 81
rect 174 80 175 81
rect 185 80 186 81
rect 186 80 187 81
rect 187 80 188 81
rect 188 80 189 81
rect 189 80 190 81
rect 190 80 191 81
rect 218 80 219 81
rect 219 80 220 81
rect 220 80 221 81
rect 221 80 222 81
rect 222 80 223 81
rect 223 80 224 81
rect 224 80 225 81
rect 225 80 226 81
rect 42 79 43 80
rect 43 79 44 80
rect 44 79 45 80
rect 45 79 46 80
rect 46 79 47 80
rect 94 79 95 80
rect 95 79 96 80
rect 96 79 97 80
rect 97 79 98 80
rect 98 79 99 80
rect 99 79 100 80
rect 100 79 101 80
rect 101 79 102 80
rect 123 79 124 80
rect 124 79 125 80
rect 125 79 126 80
rect 126 79 127 80
rect 157 79 158 80
rect 158 79 159 80
rect 159 79 160 80
rect 160 79 161 80
rect 161 79 162 80
rect 162 79 163 80
rect 163 79 164 80
rect 164 79 165 80
rect 173 79 174 80
rect 174 79 175 80
rect 185 79 186 80
rect 186 79 187 80
rect 187 79 188 80
rect 188 79 189 80
rect 189 79 190 80
rect 190 79 191 80
rect 217 79 218 80
rect 218 79 219 80
rect 219 79 220 80
rect 220 79 221 80
rect 221 79 222 80
rect 222 79 223 80
rect 223 79 224 80
rect 224 79 225 80
rect 42 78 43 79
rect 43 78 44 79
rect 44 78 45 79
rect 45 78 46 79
rect 46 78 47 79
rect 93 78 94 79
rect 94 78 95 79
rect 95 78 96 79
rect 97 78 98 79
rect 98 78 99 79
rect 99 78 100 79
rect 100 78 101 79
rect 101 78 102 79
rect 102 78 103 79
rect 123 78 124 79
rect 124 78 125 79
rect 125 78 126 79
rect 126 78 127 79
rect 158 78 159 79
rect 159 78 160 79
rect 160 78 161 79
rect 161 78 162 79
rect 162 78 163 79
rect 163 78 164 79
rect 164 78 165 79
rect 173 78 174 79
rect 174 78 175 79
rect 185 78 186 79
rect 186 78 187 79
rect 187 78 188 79
rect 188 78 189 79
rect 189 78 190 79
rect 190 78 191 79
rect 217 78 218 79
rect 218 78 219 79
rect 219 78 220 79
rect 220 78 221 79
rect 221 78 222 79
rect 222 78 223 79
rect 223 78 224 79
rect 224 78 225 79
rect 42 77 43 78
rect 43 77 44 78
rect 44 77 45 78
rect 45 77 46 78
rect 46 77 47 78
rect 92 77 93 78
rect 93 77 94 78
rect 94 77 95 78
rect 95 77 96 78
rect 97 77 98 78
rect 98 77 99 78
rect 99 77 100 78
rect 100 77 101 78
rect 101 77 102 78
rect 102 77 103 78
rect 122 77 123 78
rect 123 77 124 78
rect 124 77 125 78
rect 125 77 126 78
rect 126 77 127 78
rect 127 77 128 78
rect 159 77 160 78
rect 160 77 161 78
rect 161 77 162 78
rect 162 77 163 78
rect 163 77 164 78
rect 164 77 165 78
rect 185 77 186 78
rect 186 77 187 78
rect 187 77 188 78
rect 188 77 189 78
rect 189 77 190 78
rect 190 77 191 78
rect 217 77 218 78
rect 218 77 219 78
rect 219 77 220 78
rect 220 77 221 78
rect 221 77 222 78
rect 222 77 223 78
rect 223 77 224 78
rect 42 76 43 77
rect 43 76 44 77
rect 44 76 45 77
rect 45 76 46 77
rect 46 76 47 77
rect 92 76 93 77
rect 93 76 94 77
rect 94 76 95 77
rect 95 76 96 77
rect 97 76 98 77
rect 98 76 99 77
rect 99 76 100 77
rect 100 76 101 77
rect 101 76 102 77
rect 102 76 103 77
rect 122 76 123 77
rect 123 76 124 77
rect 124 76 125 77
rect 125 76 126 77
rect 126 76 127 77
rect 127 76 128 77
rect 140 76 141 77
rect 141 76 142 77
rect 142 76 143 77
rect 143 76 144 77
rect 144 76 145 77
rect 145 76 146 77
rect 146 76 147 77
rect 147 76 148 77
rect 148 76 149 77
rect 149 76 150 77
rect 150 76 151 77
rect 151 76 152 77
rect 159 76 160 77
rect 160 76 161 77
rect 161 76 162 77
rect 162 76 163 77
rect 163 76 164 77
rect 164 76 165 77
rect 165 76 166 77
rect 185 76 186 77
rect 186 76 187 77
rect 187 76 188 77
rect 188 76 189 77
rect 189 76 190 77
rect 190 76 191 77
rect 216 76 217 77
rect 217 76 218 77
rect 218 76 219 77
rect 219 76 220 77
rect 220 76 221 77
rect 221 76 222 77
rect 222 76 223 77
rect 223 76 224 77
rect 42 75 43 76
rect 43 75 44 76
rect 44 75 45 76
rect 45 75 46 76
rect 46 75 47 76
rect 92 75 93 76
rect 93 75 94 76
rect 94 75 95 76
rect 95 75 96 76
rect 98 75 99 76
rect 99 75 100 76
rect 100 75 101 76
rect 101 75 102 76
rect 102 75 103 76
rect 103 75 104 76
rect 122 75 123 76
rect 123 75 124 76
rect 124 75 125 76
rect 125 75 126 76
rect 126 75 127 76
rect 127 75 128 76
rect 128 75 129 76
rect 140 75 141 76
rect 141 75 142 76
rect 142 75 143 76
rect 143 75 144 76
rect 144 75 145 76
rect 145 75 146 76
rect 146 75 147 76
rect 147 75 148 76
rect 148 75 149 76
rect 149 75 150 76
rect 150 75 151 76
rect 151 75 152 76
rect 160 75 161 76
rect 161 75 162 76
rect 162 75 163 76
rect 163 75 164 76
rect 164 75 165 76
rect 165 75 166 76
rect 166 75 167 76
rect 186 75 187 76
rect 187 75 188 76
rect 188 75 189 76
rect 189 75 190 76
rect 190 75 191 76
rect 216 75 217 76
rect 217 75 218 76
rect 218 75 219 76
rect 219 75 220 76
rect 220 75 221 76
rect 221 75 222 76
rect 222 75 223 76
rect 43 74 44 75
rect 44 74 45 75
rect 45 74 46 75
rect 46 74 47 75
rect 47 74 48 75
rect 91 74 92 75
rect 92 74 93 75
rect 93 74 94 75
rect 94 74 95 75
rect 98 74 99 75
rect 99 74 100 75
rect 100 74 101 75
rect 101 74 102 75
rect 102 74 103 75
rect 103 74 104 75
rect 121 74 122 75
rect 122 74 123 75
rect 123 74 124 75
rect 124 74 125 75
rect 125 74 126 75
rect 126 74 127 75
rect 127 74 128 75
rect 128 74 129 75
rect 141 74 142 75
rect 142 74 143 75
rect 143 74 144 75
rect 144 74 145 75
rect 145 74 146 75
rect 146 74 147 75
rect 147 74 148 75
rect 148 74 149 75
rect 149 74 150 75
rect 150 74 151 75
rect 151 74 152 75
rect 160 74 161 75
rect 161 74 162 75
rect 162 74 163 75
rect 163 74 164 75
rect 164 74 165 75
rect 165 74 166 75
rect 166 74 167 75
rect 167 74 168 75
rect 185 74 186 75
rect 186 74 187 75
rect 187 74 188 75
rect 188 74 189 75
rect 189 74 190 75
rect 190 74 191 75
rect 191 74 192 75
rect 215 74 216 75
rect 216 74 217 75
rect 217 74 218 75
rect 218 74 219 75
rect 219 74 220 75
rect 220 74 221 75
rect 221 74 222 75
rect 222 74 223 75
rect 43 73 44 74
rect 44 73 45 74
rect 45 73 46 74
rect 46 73 47 74
rect 47 73 48 74
rect 48 73 49 74
rect 91 73 92 74
rect 92 73 93 74
rect 93 73 94 74
rect 94 73 95 74
rect 99 73 100 74
rect 100 73 101 74
rect 101 73 102 74
rect 102 73 103 74
rect 103 73 104 74
rect 120 73 121 74
rect 121 73 122 74
rect 122 73 123 74
rect 123 73 124 74
rect 124 73 125 74
rect 125 73 126 74
rect 126 73 127 74
rect 127 73 128 74
rect 128 73 129 74
rect 144 73 145 74
rect 145 73 146 74
rect 146 73 147 74
rect 147 73 148 74
rect 148 73 149 74
rect 161 73 162 74
rect 162 73 163 74
rect 163 73 164 74
rect 164 73 165 74
rect 165 73 166 74
rect 166 73 167 74
rect 167 73 168 74
rect 168 73 169 74
rect 182 73 183 74
rect 183 73 184 74
rect 184 73 185 74
rect 185 73 186 74
rect 186 73 187 74
rect 187 73 188 74
rect 188 73 189 74
rect 189 73 190 74
rect 190 73 191 74
rect 191 73 192 74
rect 192 73 193 74
rect 193 73 194 74
rect 194 73 195 74
rect 214 73 215 74
rect 215 73 216 74
rect 216 73 217 74
rect 217 73 218 74
rect 218 73 219 74
rect 219 73 220 74
rect 220 73 221 74
rect 221 73 222 74
rect 222 73 223 74
rect 44 72 45 73
rect 45 72 46 73
rect 46 72 47 73
rect 47 72 48 73
rect 48 72 49 73
rect 91 72 92 73
rect 92 72 93 73
rect 93 72 94 73
rect 99 72 100 73
rect 100 72 101 73
rect 101 72 102 73
rect 102 72 103 73
rect 103 72 104 73
rect 104 72 105 73
rect 120 72 121 73
rect 121 72 122 73
rect 122 72 123 73
rect 123 72 124 73
rect 124 72 125 73
rect 125 72 126 73
rect 126 72 127 73
rect 127 72 128 73
rect 128 72 129 73
rect 144 72 145 73
rect 145 72 146 73
rect 146 72 147 73
rect 147 72 148 73
rect 148 72 149 73
rect 162 72 163 73
rect 163 72 164 73
rect 164 72 165 73
rect 165 72 166 73
rect 166 72 167 73
rect 167 72 168 73
rect 168 72 169 73
rect 182 72 183 73
rect 183 72 184 73
rect 184 72 185 73
rect 185 72 186 73
rect 186 72 187 73
rect 187 72 188 73
rect 188 72 189 73
rect 189 72 190 73
rect 190 72 191 73
rect 191 72 192 73
rect 192 72 193 73
rect 193 72 194 73
rect 194 72 195 73
rect 213 72 214 73
rect 214 72 215 73
rect 215 72 216 73
rect 216 72 217 73
rect 217 72 218 73
rect 218 72 219 73
rect 219 72 220 73
rect 220 72 221 73
rect 221 72 222 73
rect 44 71 45 72
rect 45 71 46 72
rect 46 71 47 72
rect 47 71 48 72
rect 48 71 49 72
rect 49 71 50 72
rect 91 71 92 72
rect 92 71 93 72
rect 93 71 94 72
rect 99 71 100 72
rect 100 71 101 72
rect 101 71 102 72
rect 102 71 103 72
rect 103 71 104 72
rect 104 71 105 72
rect 120 71 121 72
rect 121 71 122 72
rect 122 71 123 72
rect 123 71 124 72
rect 124 71 125 72
rect 125 71 126 72
rect 126 71 127 72
rect 127 71 128 72
rect 128 71 129 72
rect 129 71 130 72
rect 144 71 145 72
rect 145 71 146 72
rect 146 71 147 72
rect 147 71 148 72
rect 148 71 149 72
rect 163 71 164 72
rect 164 71 165 72
rect 165 71 166 72
rect 166 71 167 72
rect 167 71 168 72
rect 168 71 169 72
rect 213 71 214 72
rect 214 71 215 72
rect 215 71 216 72
rect 216 71 217 72
rect 217 71 218 72
rect 218 71 219 72
rect 219 71 220 72
rect 220 71 221 72
rect 221 71 222 72
rect 45 70 46 71
rect 46 70 47 71
rect 47 70 48 71
rect 48 70 49 71
rect 49 70 50 71
rect 91 70 92 71
rect 92 70 93 71
rect 93 70 94 71
rect 99 70 100 71
rect 100 70 101 71
rect 101 70 102 71
rect 102 70 103 71
rect 103 70 104 71
rect 104 70 105 71
rect 119 70 120 71
rect 120 70 121 71
rect 121 70 122 71
rect 122 70 123 71
rect 124 70 125 71
rect 125 70 126 71
rect 126 70 127 71
rect 127 70 128 71
rect 128 70 129 71
rect 129 70 130 71
rect 144 70 145 71
rect 145 70 146 71
rect 146 70 147 71
rect 147 70 148 71
rect 148 70 149 71
rect 164 70 165 71
rect 165 70 166 71
rect 166 70 167 71
rect 167 70 168 71
rect 212 70 213 71
rect 213 70 214 71
rect 214 70 215 71
rect 215 70 216 71
rect 216 70 217 71
rect 217 70 218 71
rect 218 70 219 71
rect 219 70 220 71
rect 220 70 221 71
rect 221 70 222 71
rect 45 69 46 70
rect 46 69 47 70
rect 47 69 48 70
rect 48 69 49 70
rect 49 69 50 70
rect 50 69 51 70
rect 90 69 91 70
rect 91 69 92 70
rect 92 69 93 70
rect 100 69 101 70
rect 101 69 102 70
rect 102 69 103 70
rect 103 69 104 70
rect 104 69 105 70
rect 105 69 106 70
rect 119 69 120 70
rect 120 69 121 70
rect 121 69 122 70
rect 122 69 123 70
rect 125 69 126 70
rect 126 69 127 70
rect 127 69 128 70
rect 128 69 129 70
rect 129 69 130 70
rect 130 69 131 70
rect 144 69 145 70
rect 145 69 146 70
rect 146 69 147 70
rect 147 69 148 70
rect 148 69 149 70
rect 163 69 164 70
rect 164 69 165 70
rect 165 69 166 70
rect 166 69 167 70
rect 212 69 213 70
rect 213 69 214 70
rect 214 69 215 70
rect 215 69 216 70
rect 216 69 217 70
rect 217 69 218 70
rect 218 69 219 70
rect 219 69 220 70
rect 220 69 221 70
rect 46 68 47 69
rect 47 68 48 69
rect 48 68 49 69
rect 49 68 50 69
rect 50 68 51 69
rect 90 68 91 69
rect 91 68 92 69
rect 92 68 93 69
rect 100 68 101 69
rect 101 68 102 69
rect 102 68 103 69
rect 103 68 104 69
rect 104 68 105 69
rect 105 68 106 69
rect 119 68 120 69
rect 120 68 121 69
rect 121 68 122 69
rect 122 68 123 69
rect 125 68 126 69
rect 126 68 127 69
rect 127 68 128 69
rect 128 68 129 69
rect 129 68 130 69
rect 130 68 131 69
rect 144 68 145 69
rect 145 68 146 69
rect 146 68 147 69
rect 147 68 148 69
rect 148 68 149 69
rect 163 68 164 69
rect 164 68 165 69
rect 165 68 166 69
rect 166 68 167 69
rect 211 68 212 69
rect 212 68 213 69
rect 213 68 214 69
rect 214 68 215 69
rect 215 68 216 69
rect 216 68 217 69
rect 217 68 218 69
rect 218 68 219 69
rect 219 68 220 69
rect 220 68 221 69
rect 46 67 47 68
rect 47 67 48 68
rect 48 67 49 68
rect 49 67 50 68
rect 50 67 51 68
rect 89 67 90 68
rect 90 67 91 68
rect 91 67 92 68
rect 92 67 93 68
rect 100 67 101 68
rect 101 67 102 68
rect 102 67 103 68
rect 103 67 104 68
rect 104 67 105 68
rect 105 67 106 68
rect 106 67 107 68
rect 119 67 120 68
rect 120 67 121 68
rect 121 67 122 68
rect 125 67 126 68
rect 126 67 127 68
rect 127 67 128 68
rect 128 67 129 68
rect 129 67 130 68
rect 130 67 131 68
rect 144 67 145 68
rect 145 67 146 68
rect 146 67 147 68
rect 147 67 148 68
rect 148 67 149 68
rect 161 67 162 68
rect 162 67 163 68
rect 163 67 164 68
rect 164 67 165 68
rect 210 67 211 68
rect 211 67 212 68
rect 212 67 213 68
rect 213 67 214 68
rect 214 67 215 68
rect 215 67 216 68
rect 216 67 217 68
rect 217 67 218 68
rect 218 67 219 68
rect 219 67 220 68
rect 46 66 47 67
rect 47 66 48 67
rect 48 66 49 67
rect 49 66 50 67
rect 50 66 51 67
rect 51 66 52 67
rect 89 66 90 67
rect 90 66 91 67
rect 91 66 92 67
rect 101 66 102 67
rect 102 66 103 67
rect 103 66 104 67
rect 104 66 105 67
rect 105 66 106 67
rect 106 66 107 67
rect 118 66 119 67
rect 119 66 120 67
rect 120 66 121 67
rect 121 66 122 67
rect 126 66 127 67
rect 127 66 128 67
rect 128 66 129 67
rect 129 66 130 67
rect 130 66 131 67
rect 131 66 132 67
rect 144 66 145 67
rect 145 66 146 67
rect 146 66 147 67
rect 147 66 148 67
rect 148 66 149 67
rect 160 66 161 67
rect 161 66 162 67
rect 162 66 163 67
rect 163 66 164 67
rect 164 66 165 67
rect 209 66 210 67
rect 210 66 211 67
rect 211 66 212 67
rect 212 66 213 67
rect 213 66 214 67
rect 214 66 215 67
rect 215 66 216 67
rect 216 66 217 67
rect 217 66 218 67
rect 218 66 219 67
rect 219 66 220 67
rect 46 65 47 66
rect 47 65 48 66
rect 48 65 49 66
rect 49 65 50 66
rect 50 65 51 66
rect 51 65 52 66
rect 88 65 89 66
rect 89 65 90 66
rect 90 65 91 66
rect 91 65 92 66
rect 102 65 103 66
rect 103 65 104 66
rect 104 65 105 66
rect 105 65 106 66
rect 106 65 107 66
rect 107 65 108 66
rect 118 65 119 66
rect 119 65 120 66
rect 120 65 121 66
rect 127 65 128 66
rect 128 65 129 66
rect 129 65 130 66
rect 130 65 131 66
rect 131 65 132 66
rect 132 65 133 66
rect 144 65 145 66
rect 145 65 146 66
rect 146 65 147 66
rect 147 65 148 66
rect 148 65 149 66
rect 160 65 161 66
rect 161 65 162 66
rect 162 65 163 66
rect 163 65 164 66
rect 175 65 176 66
rect 176 65 177 66
rect 209 65 210 66
rect 210 65 211 66
rect 211 65 212 66
rect 212 65 213 66
rect 213 65 214 66
rect 214 65 215 66
rect 215 65 216 66
rect 216 65 217 66
rect 217 65 218 66
rect 47 64 48 65
rect 48 64 49 65
rect 49 64 50 65
rect 50 64 51 65
rect 51 64 52 65
rect 52 64 53 65
rect 88 64 89 65
rect 89 64 90 65
rect 90 64 91 65
rect 91 64 92 65
rect 102 64 103 65
rect 103 64 104 65
rect 104 64 105 65
rect 105 64 106 65
rect 106 64 107 65
rect 107 64 108 65
rect 118 64 119 65
rect 119 64 120 65
rect 120 64 121 65
rect 127 64 128 65
rect 128 64 129 65
rect 129 64 130 65
rect 130 64 131 65
rect 131 64 132 65
rect 132 64 133 65
rect 144 64 145 65
rect 145 64 146 65
rect 146 64 147 65
rect 147 64 148 65
rect 148 64 149 65
rect 159 64 160 65
rect 160 64 161 65
rect 161 64 162 65
rect 162 64 163 65
rect 163 64 164 65
rect 174 64 175 65
rect 175 64 176 65
rect 176 64 177 65
rect 208 64 209 65
rect 209 64 210 65
rect 210 64 211 65
rect 211 64 212 65
rect 212 64 213 65
rect 213 64 214 65
rect 214 64 215 65
rect 215 64 216 65
rect 216 64 217 65
rect 217 64 218 65
rect 47 63 48 64
rect 48 63 49 64
rect 49 63 50 64
rect 50 63 51 64
rect 51 63 52 64
rect 52 63 53 64
rect 88 63 89 64
rect 89 63 90 64
rect 90 63 91 64
rect 91 63 92 64
rect 102 63 103 64
rect 103 63 104 64
rect 104 63 105 64
rect 105 63 106 64
rect 106 63 107 64
rect 107 63 108 64
rect 117 63 118 64
rect 118 63 119 64
rect 119 63 120 64
rect 127 63 128 64
rect 128 63 129 64
rect 129 63 130 64
rect 130 63 131 64
rect 131 63 132 64
rect 132 63 133 64
rect 144 63 145 64
rect 145 63 146 64
rect 146 63 147 64
rect 147 63 148 64
rect 148 63 149 64
rect 158 63 159 64
rect 159 63 160 64
rect 160 63 161 64
rect 161 63 162 64
rect 174 63 175 64
rect 175 63 176 64
rect 176 63 177 64
rect 207 63 208 64
rect 208 63 209 64
rect 209 63 210 64
rect 210 63 211 64
rect 211 63 212 64
rect 212 63 213 64
rect 213 63 214 64
rect 214 63 215 64
rect 215 63 216 64
rect 216 63 217 64
rect 48 62 49 63
rect 49 62 50 63
rect 50 62 51 63
rect 51 62 52 63
rect 52 62 53 63
rect 53 62 54 63
rect 87 62 88 63
rect 88 62 89 63
rect 89 62 90 63
rect 90 62 91 63
rect 91 62 92 63
rect 102 62 103 63
rect 103 62 104 63
rect 104 62 105 63
rect 105 62 106 63
rect 106 62 107 63
rect 107 62 108 63
rect 108 62 109 63
rect 117 62 118 63
rect 118 62 119 63
rect 119 62 120 63
rect 128 62 129 63
rect 129 62 130 63
rect 130 62 131 63
rect 131 62 132 63
rect 132 62 133 63
rect 144 62 145 63
rect 145 62 146 63
rect 146 62 147 63
rect 147 62 148 63
rect 148 62 149 63
rect 158 62 159 63
rect 159 62 160 63
rect 160 62 161 63
rect 161 62 162 63
rect 173 62 174 63
rect 174 62 175 63
rect 175 62 176 63
rect 176 62 177 63
rect 206 62 207 63
rect 207 62 208 63
rect 208 62 209 63
rect 209 62 210 63
rect 210 62 211 63
rect 211 62 212 63
rect 212 62 213 63
rect 213 62 214 63
rect 214 62 215 63
rect 215 62 216 63
rect 48 61 49 62
rect 49 61 50 62
rect 50 61 51 62
rect 51 61 52 62
rect 52 61 53 62
rect 53 61 54 62
rect 54 61 55 62
rect 85 61 86 62
rect 86 61 87 62
rect 87 61 88 62
rect 88 61 89 62
rect 89 61 90 62
rect 90 61 91 62
rect 91 61 92 62
rect 101 61 102 62
rect 102 61 103 62
rect 103 61 104 62
rect 104 61 105 62
rect 105 61 106 62
rect 106 61 107 62
rect 107 61 108 62
rect 108 61 109 62
rect 109 61 110 62
rect 117 61 118 62
rect 118 61 119 62
rect 119 61 120 62
rect 128 61 129 62
rect 129 61 130 62
rect 130 61 131 62
rect 131 61 132 62
rect 132 61 133 62
rect 144 61 145 62
rect 145 61 146 62
rect 146 61 147 62
rect 147 61 148 62
rect 148 61 149 62
rect 156 61 157 62
rect 157 61 158 62
rect 158 61 159 62
rect 159 61 160 62
rect 160 61 161 62
rect 172 61 173 62
rect 173 61 174 62
rect 174 61 175 62
rect 175 61 176 62
rect 176 61 177 62
rect 205 61 206 62
rect 206 61 207 62
rect 207 61 208 62
rect 208 61 209 62
rect 209 61 210 62
rect 210 61 211 62
rect 211 61 212 62
rect 212 61 213 62
rect 213 61 214 62
rect 214 61 215 62
rect 49 60 50 61
rect 50 60 51 61
rect 51 60 52 61
rect 52 60 53 61
rect 53 60 54 61
rect 54 60 55 61
rect 84 60 85 61
rect 85 60 86 61
rect 86 60 87 61
rect 87 60 88 61
rect 88 60 89 61
rect 89 60 90 61
rect 90 60 91 61
rect 91 60 92 61
rect 92 60 93 61
rect 93 60 94 61
rect 99 60 100 61
rect 100 60 101 61
rect 101 60 102 61
rect 102 60 103 61
rect 103 60 104 61
rect 104 60 105 61
rect 105 60 106 61
rect 106 60 107 61
rect 107 60 108 61
rect 108 60 109 61
rect 109 60 110 61
rect 110 60 111 61
rect 111 60 112 61
rect 116 60 117 61
rect 117 60 118 61
rect 118 60 119 61
rect 119 60 120 61
rect 128 60 129 61
rect 129 60 130 61
rect 130 60 131 61
rect 131 60 132 61
rect 132 60 133 61
rect 133 60 134 61
rect 144 60 145 61
rect 145 60 146 61
rect 146 60 147 61
rect 147 60 148 61
rect 148 60 149 61
rect 156 60 157 61
rect 157 60 158 61
rect 158 60 159 61
rect 159 60 160 61
rect 160 60 161 61
rect 161 60 162 61
rect 162 60 163 61
rect 163 60 164 61
rect 164 60 165 61
rect 165 60 166 61
rect 166 60 167 61
rect 167 60 168 61
rect 168 60 169 61
rect 169 60 170 61
rect 170 60 171 61
rect 171 60 172 61
rect 172 60 173 61
rect 173 60 174 61
rect 174 60 175 61
rect 175 60 176 61
rect 176 60 177 61
rect 205 60 206 61
rect 206 60 207 61
rect 207 60 208 61
rect 208 60 209 61
rect 209 60 210 61
rect 210 60 211 61
rect 211 60 212 61
rect 212 60 213 61
rect 213 60 214 61
rect 214 60 215 61
rect 49 59 50 60
rect 50 59 51 60
rect 51 59 52 60
rect 52 59 53 60
rect 53 59 54 60
rect 54 59 55 60
rect 55 59 56 60
rect 84 59 85 60
rect 85 59 86 60
rect 86 59 87 60
rect 87 59 88 60
rect 88 59 89 60
rect 89 59 90 60
rect 90 59 91 60
rect 91 59 92 60
rect 92 59 93 60
rect 93 59 94 60
rect 99 59 100 60
rect 100 59 101 60
rect 101 59 102 60
rect 102 59 103 60
rect 103 59 104 60
rect 104 59 105 60
rect 105 59 106 60
rect 106 59 107 60
rect 107 59 108 60
rect 108 59 109 60
rect 109 59 110 60
rect 110 59 111 60
rect 111 59 112 60
rect 116 59 117 60
rect 117 59 118 60
rect 118 59 119 60
rect 119 59 120 60
rect 128 59 129 60
rect 129 59 130 60
rect 130 59 131 60
rect 131 59 132 60
rect 132 59 133 60
rect 133 59 134 60
rect 134 59 135 60
rect 144 59 145 60
rect 145 59 146 60
rect 146 59 147 60
rect 147 59 148 60
rect 148 59 149 60
rect 155 59 156 60
rect 156 59 157 60
rect 157 59 158 60
rect 158 59 159 60
rect 159 59 160 60
rect 160 59 161 60
rect 161 59 162 60
rect 162 59 163 60
rect 163 59 164 60
rect 164 59 165 60
rect 165 59 166 60
rect 166 59 167 60
rect 167 59 168 60
rect 168 59 169 60
rect 169 59 170 60
rect 170 59 171 60
rect 171 59 172 60
rect 172 59 173 60
rect 173 59 174 60
rect 174 59 175 60
rect 175 59 176 60
rect 203 59 204 60
rect 204 59 205 60
rect 205 59 206 60
rect 206 59 207 60
rect 207 59 208 60
rect 208 59 209 60
rect 209 59 210 60
rect 210 59 211 60
rect 211 59 212 60
rect 212 59 213 60
rect 213 59 214 60
rect 50 58 51 59
rect 51 58 52 59
rect 52 58 53 59
rect 53 58 54 59
rect 54 58 55 59
rect 55 58 56 59
rect 115 58 116 59
rect 116 58 117 59
rect 117 58 118 59
rect 118 58 119 59
rect 129 58 130 59
rect 130 58 131 59
rect 131 58 132 59
rect 132 58 133 59
rect 133 58 134 59
rect 134 58 135 59
rect 144 58 145 59
rect 145 58 146 59
rect 146 58 147 59
rect 147 58 148 59
rect 148 58 149 59
rect 154 58 155 59
rect 155 58 156 59
rect 156 58 157 59
rect 157 58 158 59
rect 158 58 159 59
rect 159 58 160 59
rect 160 58 161 59
rect 161 58 162 59
rect 162 58 163 59
rect 163 58 164 59
rect 164 58 165 59
rect 165 58 166 59
rect 166 58 167 59
rect 167 58 168 59
rect 168 58 169 59
rect 169 58 170 59
rect 170 58 171 59
rect 171 58 172 59
rect 172 58 173 59
rect 173 58 174 59
rect 174 58 175 59
rect 175 58 176 59
rect 202 58 203 59
rect 203 58 204 59
rect 204 58 205 59
rect 205 58 206 59
rect 206 58 207 59
rect 207 58 208 59
rect 208 58 209 59
rect 209 58 210 59
rect 210 58 211 59
rect 211 58 212 59
rect 212 58 213 59
rect 50 57 51 58
rect 51 57 52 58
rect 52 57 53 58
rect 53 57 54 58
rect 54 57 55 58
rect 55 57 56 58
rect 56 57 57 58
rect 115 57 116 58
rect 116 57 117 58
rect 117 57 118 58
rect 118 57 119 58
rect 129 57 130 58
rect 130 57 131 58
rect 131 57 132 58
rect 132 57 133 58
rect 133 57 134 58
rect 134 57 135 58
rect 135 57 136 58
rect 144 57 145 58
rect 145 57 146 58
rect 146 57 147 58
rect 147 57 148 58
rect 148 57 149 58
rect 153 57 154 58
rect 154 57 155 58
rect 155 57 156 58
rect 156 57 157 58
rect 157 57 158 58
rect 158 57 159 58
rect 159 57 160 58
rect 160 57 161 58
rect 161 57 162 58
rect 162 57 163 58
rect 163 57 164 58
rect 164 57 165 58
rect 165 57 166 58
rect 166 57 167 58
rect 167 57 168 58
rect 168 57 169 58
rect 169 57 170 58
rect 170 57 171 58
rect 171 57 172 58
rect 172 57 173 58
rect 173 57 174 58
rect 174 57 175 58
rect 175 57 176 58
rect 201 57 202 58
rect 202 57 203 58
rect 203 57 204 58
rect 204 57 205 58
rect 205 57 206 58
rect 206 57 207 58
rect 207 57 208 58
rect 208 57 209 58
rect 209 57 210 58
rect 210 57 211 58
rect 51 56 52 57
rect 52 56 53 57
rect 53 56 54 57
rect 54 56 55 57
rect 55 56 56 57
rect 56 56 57 57
rect 57 56 58 57
rect 115 56 116 57
rect 116 56 117 57
rect 117 56 118 57
rect 118 56 119 57
rect 129 56 130 57
rect 130 56 131 57
rect 131 56 132 57
rect 132 56 133 57
rect 133 56 134 57
rect 134 56 135 57
rect 135 56 136 57
rect 144 56 145 57
rect 145 56 146 57
rect 146 56 147 57
rect 147 56 148 57
rect 148 56 149 57
rect 153 56 154 57
rect 154 56 155 57
rect 155 56 156 57
rect 156 56 157 57
rect 157 56 158 57
rect 158 56 159 57
rect 159 56 160 57
rect 160 56 161 57
rect 161 56 162 57
rect 162 56 163 57
rect 163 56 164 57
rect 164 56 165 57
rect 165 56 166 57
rect 166 56 167 57
rect 167 56 168 57
rect 168 56 169 57
rect 169 56 170 57
rect 170 56 171 57
rect 171 56 172 57
rect 172 56 173 57
rect 173 56 174 57
rect 174 56 175 57
rect 201 56 202 57
rect 202 56 203 57
rect 203 56 204 57
rect 204 56 205 57
rect 205 56 206 57
rect 206 56 207 57
rect 207 56 208 57
rect 208 56 209 57
rect 209 56 210 57
rect 210 56 211 57
rect 51 55 52 56
rect 52 55 53 56
rect 53 55 54 56
rect 54 55 55 56
rect 55 55 56 56
rect 56 55 57 56
rect 57 55 58 56
rect 113 55 114 56
rect 114 55 115 56
rect 115 55 116 56
rect 116 55 117 56
rect 117 55 118 56
rect 118 55 119 56
rect 129 55 130 56
rect 130 55 131 56
rect 131 55 132 56
rect 132 55 133 56
rect 133 55 134 56
rect 134 55 135 56
rect 135 55 136 56
rect 136 55 137 56
rect 144 55 145 56
rect 145 55 146 56
rect 146 55 147 56
rect 147 55 148 56
rect 148 55 149 56
rect 199 55 200 56
rect 200 55 201 56
rect 201 55 202 56
rect 202 55 203 56
rect 203 55 204 56
rect 204 55 205 56
rect 205 55 206 56
rect 206 55 207 56
rect 207 55 208 56
rect 208 55 209 56
rect 209 55 210 56
rect 52 54 53 55
rect 53 54 54 55
rect 54 54 55 55
rect 55 54 56 55
rect 56 54 57 55
rect 57 54 58 55
rect 58 54 59 55
rect 111 54 112 55
rect 112 54 113 55
rect 113 54 114 55
rect 114 54 115 55
rect 115 54 116 55
rect 116 54 117 55
rect 117 54 118 55
rect 118 54 119 55
rect 119 54 120 55
rect 120 54 121 55
rect 127 54 128 55
rect 128 54 129 55
rect 129 54 130 55
rect 130 54 131 55
rect 131 54 132 55
rect 132 54 133 55
rect 133 54 134 55
rect 134 54 135 55
rect 135 54 136 55
rect 136 54 137 55
rect 137 54 138 55
rect 138 54 139 55
rect 144 54 145 55
rect 145 54 146 55
rect 146 54 147 55
rect 147 54 148 55
rect 148 54 149 55
rect 198 54 199 55
rect 199 54 200 55
rect 200 54 201 55
rect 201 54 202 55
rect 202 54 203 55
rect 203 54 204 55
rect 204 54 205 55
rect 205 54 206 55
rect 206 54 207 55
rect 207 54 208 55
rect 208 54 209 55
rect 209 54 210 55
rect 53 53 54 54
rect 54 53 55 54
rect 55 53 56 54
rect 56 53 57 54
rect 57 53 58 54
rect 58 53 59 54
rect 111 53 112 54
rect 112 53 113 54
rect 113 53 114 54
rect 114 53 115 54
rect 115 53 116 54
rect 116 53 117 54
rect 117 53 118 54
rect 118 53 119 54
rect 119 53 120 54
rect 120 53 121 54
rect 127 53 128 54
rect 128 53 129 54
rect 129 53 130 54
rect 130 53 131 54
rect 131 53 132 54
rect 132 53 133 54
rect 133 53 134 54
rect 134 53 135 54
rect 135 53 136 54
rect 136 53 137 54
rect 137 53 138 54
rect 138 53 139 54
rect 144 53 145 54
rect 145 53 146 54
rect 146 53 147 54
rect 147 53 148 54
rect 148 53 149 54
rect 197 53 198 54
rect 198 53 199 54
rect 199 53 200 54
rect 200 53 201 54
rect 201 53 202 54
rect 202 53 203 54
rect 203 53 204 54
rect 204 53 205 54
rect 205 53 206 54
rect 206 53 207 54
rect 207 53 208 54
rect 208 53 209 54
rect 53 52 54 53
rect 54 52 55 53
rect 55 52 56 53
rect 56 52 57 53
rect 57 52 58 53
rect 58 52 59 53
rect 59 52 60 53
rect 113 52 114 53
rect 114 52 115 53
rect 115 52 116 53
rect 116 52 117 53
rect 118 52 119 53
rect 119 52 120 53
rect 128 52 129 53
rect 129 52 130 53
rect 130 52 131 53
rect 131 52 132 53
rect 133 52 134 53
rect 134 52 135 53
rect 135 52 136 53
rect 144 52 145 53
rect 145 52 146 53
rect 146 52 147 53
rect 147 52 148 53
rect 148 52 149 53
rect 195 52 196 53
rect 196 52 197 53
rect 197 52 198 53
rect 198 52 199 53
rect 199 52 200 53
rect 200 52 201 53
rect 201 52 202 53
rect 202 52 203 53
rect 203 52 204 53
rect 204 52 205 53
rect 205 52 206 53
rect 206 52 207 53
rect 54 51 55 52
rect 55 51 56 52
rect 56 51 57 52
rect 57 51 58 52
rect 58 51 59 52
rect 59 51 60 52
rect 60 51 61 52
rect 144 51 145 52
rect 145 51 146 52
rect 146 51 147 52
rect 147 51 148 52
rect 148 51 149 52
rect 194 51 195 52
rect 195 51 196 52
rect 196 51 197 52
rect 197 51 198 52
rect 198 51 199 52
rect 199 51 200 52
rect 200 51 201 52
rect 201 51 202 52
rect 202 51 203 52
rect 203 51 204 52
rect 204 51 205 52
rect 205 51 206 52
rect 54 50 55 51
rect 55 50 56 51
rect 56 50 57 51
rect 57 50 58 51
rect 58 50 59 51
rect 59 50 60 51
rect 60 50 61 51
rect 61 50 62 51
rect 144 50 145 51
rect 145 50 146 51
rect 146 50 147 51
rect 147 50 148 51
rect 148 50 149 51
rect 193 50 194 51
rect 194 50 195 51
rect 195 50 196 51
rect 196 50 197 51
rect 197 50 198 51
rect 198 50 199 51
rect 199 50 200 51
rect 200 50 201 51
rect 201 50 202 51
rect 202 50 203 51
rect 203 50 204 51
rect 204 50 205 51
rect 55 49 56 50
rect 56 49 57 50
rect 57 49 58 50
rect 58 49 59 50
rect 59 49 60 50
rect 60 49 61 50
rect 61 49 62 50
rect 62 49 63 50
rect 142 49 143 50
rect 143 49 144 50
rect 144 49 145 50
rect 145 49 146 50
rect 146 49 147 50
rect 147 49 148 50
rect 148 49 149 50
rect 149 49 150 50
rect 192 49 193 50
rect 193 49 194 50
rect 194 49 195 50
rect 195 49 196 50
rect 196 49 197 50
rect 197 49 198 50
rect 198 49 199 50
rect 199 49 200 50
rect 200 49 201 50
rect 201 49 202 50
rect 202 49 203 50
rect 203 49 204 50
rect 56 48 57 49
rect 57 48 58 49
rect 58 48 59 49
rect 59 48 60 49
rect 60 48 61 49
rect 61 48 62 49
rect 62 48 63 49
rect 63 48 64 49
rect 140 48 141 49
rect 141 48 142 49
rect 142 48 143 49
rect 143 48 144 49
rect 144 48 145 49
rect 145 48 146 49
rect 146 48 147 49
rect 147 48 148 49
rect 148 48 149 49
rect 149 48 150 49
rect 150 48 151 49
rect 151 48 152 49
rect 191 48 192 49
rect 192 48 193 49
rect 193 48 194 49
rect 194 48 195 49
rect 195 48 196 49
rect 196 48 197 49
rect 197 48 198 49
rect 198 48 199 49
rect 199 48 200 49
rect 200 48 201 49
rect 201 48 202 49
rect 202 48 203 49
rect 56 47 57 48
rect 57 47 58 48
rect 58 47 59 48
rect 59 47 60 48
rect 60 47 61 48
rect 61 47 62 48
rect 62 47 63 48
rect 63 47 64 48
rect 140 47 141 48
rect 141 47 142 48
rect 142 47 143 48
rect 143 47 144 48
rect 144 47 145 48
rect 145 47 146 48
rect 146 47 147 48
rect 147 47 148 48
rect 148 47 149 48
rect 149 47 150 48
rect 150 47 151 48
rect 151 47 152 48
rect 190 47 191 48
rect 191 47 192 48
rect 192 47 193 48
rect 193 47 194 48
rect 194 47 195 48
rect 195 47 196 48
rect 196 47 197 48
rect 197 47 198 48
rect 198 47 199 48
rect 199 47 200 48
rect 200 47 201 48
rect 201 47 202 48
rect 57 46 58 47
rect 58 46 59 47
rect 59 46 60 47
rect 60 46 61 47
rect 61 46 62 47
rect 62 46 63 47
rect 63 46 64 47
rect 189 46 190 47
rect 190 46 191 47
rect 191 46 192 47
rect 192 46 193 47
rect 193 46 194 47
rect 194 46 195 47
rect 195 46 196 47
rect 196 46 197 47
rect 197 46 198 47
rect 198 46 199 47
rect 199 46 200 47
rect 200 46 201 47
rect 58 45 59 46
rect 59 45 60 46
rect 60 45 61 46
rect 61 45 62 46
rect 62 45 63 46
rect 63 45 64 46
rect 64 45 65 46
rect 65 45 66 46
rect 187 45 188 46
rect 188 45 189 46
rect 189 45 190 46
rect 190 45 191 46
rect 191 45 192 46
rect 192 45 193 46
rect 193 45 194 46
rect 194 45 195 46
rect 195 45 196 46
rect 196 45 197 46
rect 197 45 198 46
rect 198 45 199 46
rect 199 45 200 46
rect 59 44 60 45
rect 60 44 61 45
rect 61 44 62 45
rect 62 44 63 45
rect 63 44 64 45
rect 64 44 65 45
rect 65 44 66 45
rect 66 44 67 45
rect 187 44 188 45
rect 188 44 189 45
rect 189 44 190 45
rect 190 44 191 45
rect 191 44 192 45
rect 192 44 193 45
rect 193 44 194 45
rect 194 44 195 45
rect 195 44 196 45
rect 196 44 197 45
rect 197 44 198 45
rect 59 43 60 44
rect 60 43 61 44
rect 61 43 62 44
rect 62 43 63 44
rect 63 43 64 44
rect 64 43 65 44
rect 65 43 66 44
rect 66 43 67 44
rect 67 43 68 44
rect 185 43 186 44
rect 186 43 187 44
rect 187 43 188 44
rect 188 43 189 44
rect 189 43 190 44
rect 190 43 191 44
rect 191 43 192 44
rect 192 43 193 44
rect 193 43 194 44
rect 194 43 195 44
rect 195 43 196 44
rect 196 43 197 44
rect 60 42 61 43
rect 61 42 62 43
rect 62 42 63 43
rect 63 42 64 43
rect 64 42 65 43
rect 65 42 66 43
rect 66 42 67 43
rect 67 42 68 43
rect 185 42 186 43
rect 186 42 187 43
rect 187 42 188 43
rect 188 42 189 43
rect 189 42 190 43
rect 190 42 191 43
rect 191 42 192 43
rect 192 42 193 43
rect 193 42 194 43
rect 194 42 195 43
rect 195 42 196 43
rect 61 41 62 42
rect 62 41 63 42
rect 63 41 64 42
rect 64 41 65 42
rect 65 41 66 42
rect 66 41 67 42
rect 67 41 68 42
rect 68 41 69 42
rect 69 41 70 42
rect 184 41 185 42
rect 185 41 186 42
rect 186 41 187 42
rect 187 41 188 42
rect 188 41 189 42
rect 189 41 190 42
rect 190 41 191 42
rect 191 41 192 42
rect 192 41 193 42
rect 193 41 194 42
rect 194 41 195 42
rect 62 40 63 41
rect 63 40 64 41
rect 64 40 65 41
rect 65 40 66 41
rect 66 40 67 41
rect 67 40 68 41
rect 68 40 69 41
rect 69 40 70 41
rect 183 40 184 41
rect 184 40 185 41
rect 185 40 186 41
rect 186 40 187 41
rect 187 40 188 41
rect 188 40 189 41
rect 189 40 190 41
rect 190 40 191 41
rect 191 40 192 41
rect 192 40 193 41
rect 193 40 194 41
rect 63 39 64 40
rect 64 39 65 40
rect 65 39 66 40
rect 66 39 67 40
rect 67 39 68 40
rect 68 39 69 40
rect 69 39 70 40
rect 70 39 71 40
rect 71 39 72 40
rect 181 39 182 40
rect 182 39 183 40
rect 183 39 184 40
rect 184 39 185 40
rect 185 39 186 40
rect 186 39 187 40
rect 187 39 188 40
rect 188 39 189 40
rect 189 39 190 40
rect 190 39 191 40
rect 191 39 192 40
rect 192 39 193 40
rect 64 38 65 39
rect 65 38 66 39
rect 66 38 67 39
rect 67 38 68 39
rect 68 38 69 39
rect 69 38 70 39
rect 70 38 71 39
rect 71 38 72 39
rect 72 38 73 39
rect 181 38 182 39
rect 182 38 183 39
rect 183 38 184 39
rect 184 38 185 39
rect 185 38 186 39
rect 186 38 187 39
rect 187 38 188 39
rect 188 38 189 39
rect 189 38 190 39
rect 65 37 66 38
rect 66 37 67 38
rect 67 37 68 38
rect 68 37 69 38
rect 69 37 70 38
rect 70 37 71 38
rect 71 37 72 38
rect 72 37 73 38
rect 73 37 74 38
rect 180 37 181 38
rect 181 37 182 38
rect 182 37 183 38
rect 183 37 184 38
rect 184 37 185 38
rect 185 37 186 38
rect 186 37 187 38
rect 187 37 188 38
rect 188 37 189 38
rect 189 37 190 38
rect 66 36 67 37
rect 67 36 68 37
rect 68 36 69 37
rect 69 36 70 37
rect 70 36 71 37
rect 71 36 72 37
rect 72 36 73 37
rect 73 36 74 37
rect 74 36 75 37
rect 179 36 180 37
rect 180 36 181 37
rect 181 36 182 37
rect 182 36 183 37
rect 183 36 184 37
rect 184 36 185 37
rect 185 36 186 37
rect 186 36 187 37
rect 187 36 188 37
rect 188 36 189 37
rect 67 35 68 36
rect 68 35 69 36
rect 69 35 70 36
rect 70 35 71 36
rect 71 35 72 36
rect 72 35 73 36
rect 73 35 74 36
rect 74 35 75 36
rect 75 35 76 36
rect 178 35 179 36
rect 179 35 180 36
rect 180 35 181 36
rect 181 35 182 36
rect 182 35 183 36
rect 183 35 184 36
rect 184 35 185 36
rect 185 35 186 36
rect 186 35 187 36
rect 67 34 68 35
rect 68 34 69 35
rect 69 34 70 35
rect 70 34 71 35
rect 71 34 72 35
rect 72 34 73 35
rect 73 34 74 35
rect 74 34 75 35
rect 75 34 76 35
rect 76 34 77 35
rect 177 34 178 35
rect 178 34 179 35
rect 179 34 180 35
rect 180 34 181 35
rect 181 34 182 35
rect 182 34 183 35
rect 183 34 184 35
rect 184 34 185 35
rect 185 34 186 35
rect 69 33 70 34
rect 70 33 71 34
rect 71 33 72 34
rect 72 33 73 34
rect 73 33 74 34
rect 74 33 75 34
rect 75 33 76 34
rect 76 33 77 34
rect 77 33 78 34
rect 176 33 177 34
rect 177 33 178 34
rect 178 33 179 34
rect 179 33 180 34
rect 180 33 181 34
rect 181 33 182 34
rect 182 33 183 34
rect 183 33 184 34
rect 184 33 185 34
rect 69 32 70 33
rect 70 32 71 33
rect 71 32 72 33
rect 72 32 73 33
rect 73 32 74 33
rect 74 32 75 33
rect 75 32 76 33
rect 76 32 77 33
rect 77 32 78 33
rect 78 32 79 33
rect 79 32 80 33
rect 174 32 175 33
rect 175 32 176 33
rect 176 32 177 33
rect 177 32 178 33
rect 178 32 179 33
rect 179 32 180 33
rect 180 32 181 33
rect 181 32 182 33
rect 182 32 183 33
rect 183 32 184 33
rect 71 31 72 32
rect 72 31 73 32
rect 73 31 74 32
rect 74 31 75 32
rect 75 31 76 32
rect 76 31 77 32
rect 77 31 78 32
rect 78 31 79 32
rect 79 31 80 32
rect 80 31 81 32
rect 173 31 174 32
rect 174 31 175 32
rect 175 31 176 32
rect 176 31 177 32
rect 177 31 178 32
rect 178 31 179 32
rect 179 31 180 32
rect 180 31 181 32
rect 181 31 182 32
rect 72 30 73 31
rect 73 30 74 31
rect 74 30 75 31
rect 75 30 76 31
rect 76 30 77 31
rect 77 30 78 31
rect 78 30 79 31
rect 79 30 80 31
rect 80 30 81 31
rect 81 30 82 31
rect 82 30 83 31
rect 172 30 173 31
rect 173 30 174 31
rect 174 30 175 31
rect 175 30 176 31
rect 176 30 177 31
rect 177 30 178 31
rect 178 30 179 31
rect 179 30 180 31
rect 73 29 74 30
rect 74 29 75 30
rect 75 29 76 30
rect 76 29 77 30
rect 77 29 78 30
rect 78 29 79 30
rect 79 29 80 30
rect 80 29 81 30
rect 81 29 82 30
rect 82 29 83 30
rect 83 29 84 30
rect 172 29 173 30
rect 173 29 174 30
rect 174 29 175 30
rect 175 29 176 30
rect 176 29 177 30
rect 177 29 178 30
rect 178 29 179 30
rect 75 28 76 29
rect 76 28 77 29
rect 77 28 78 29
rect 78 28 79 29
rect 79 28 80 29
rect 80 28 81 29
rect 81 28 82 29
rect 82 28 83 29
rect 83 28 84 29
rect 84 28 85 29
rect 170 28 171 29
rect 171 28 172 29
rect 172 28 173 29
rect 173 28 174 29
rect 174 28 175 29
rect 175 28 176 29
rect 176 28 177 29
rect 75 27 76 28
rect 76 27 77 28
rect 77 27 78 28
rect 78 27 79 28
rect 79 27 80 28
rect 80 27 81 28
rect 81 27 82 28
rect 82 27 83 28
rect 83 27 84 28
rect 84 27 85 28
rect 85 27 86 28
rect 86 27 87 28
rect 169 27 170 28
rect 170 27 171 28
rect 171 27 172 28
rect 172 27 173 28
rect 173 27 174 28
rect 174 27 175 28
rect 175 27 176 28
rect 176 27 177 28
rect 77 26 78 27
rect 78 26 79 27
rect 79 26 80 27
rect 80 26 81 27
rect 81 26 82 27
rect 82 26 83 27
rect 83 26 84 27
rect 84 26 85 27
rect 85 26 86 27
rect 86 26 87 27
rect 87 26 88 27
rect 136 26 137 27
rect 137 26 138 27
rect 138 26 139 27
rect 168 26 169 27
rect 169 26 170 27
rect 170 26 171 27
rect 171 26 172 27
rect 172 26 173 27
rect 173 26 174 27
rect 174 26 175 27
rect 78 25 79 26
rect 79 25 80 26
rect 80 25 81 26
rect 81 25 82 26
rect 82 25 83 26
rect 83 25 84 26
rect 84 25 85 26
rect 85 25 86 26
rect 86 25 87 26
rect 87 25 88 26
rect 88 25 89 26
rect 89 25 90 26
rect 90 25 91 26
rect 91 25 92 26
rect 92 25 93 26
rect 93 25 94 26
rect 94 25 95 26
rect 95 25 96 26
rect 96 25 97 26
rect 128 25 129 26
rect 129 25 130 26
rect 130 25 131 26
rect 131 25 132 26
rect 132 25 133 26
rect 133 25 134 26
rect 134 25 135 26
rect 135 25 136 26
rect 136 25 137 26
rect 137 25 138 26
rect 138 25 139 26
rect 166 25 167 26
rect 167 25 168 26
rect 168 25 169 26
rect 169 25 170 26
rect 170 25 171 26
rect 171 25 172 26
rect 172 25 173 26
rect 173 25 174 26
rect 80 24 81 25
rect 81 24 82 25
rect 82 24 83 25
rect 83 24 84 25
rect 84 24 85 25
rect 85 24 86 25
rect 86 24 87 25
rect 87 24 88 25
rect 88 24 89 25
rect 89 24 90 25
rect 90 24 91 25
rect 91 24 92 25
rect 92 24 93 25
rect 93 24 94 25
rect 94 24 95 25
rect 95 24 96 25
rect 96 24 97 25
rect 97 24 98 25
rect 98 24 99 25
rect 99 24 100 25
rect 100 24 101 25
rect 101 24 102 25
rect 102 24 103 25
rect 103 24 104 25
rect 104 24 105 25
rect 105 24 106 25
rect 106 24 107 25
rect 107 24 108 25
rect 119 24 120 25
rect 120 24 121 25
rect 122 24 123 25
rect 123 24 124 25
rect 124 24 125 25
rect 125 24 126 25
rect 126 24 127 25
rect 127 24 128 25
rect 128 24 129 25
rect 129 24 130 25
rect 130 24 131 25
rect 131 24 132 25
rect 132 24 133 25
rect 133 24 134 25
rect 134 24 135 25
rect 135 24 136 25
rect 136 24 137 25
rect 165 24 166 25
rect 166 24 167 25
rect 167 24 168 25
rect 168 24 169 25
rect 169 24 170 25
rect 170 24 171 25
rect 171 24 172 25
rect 82 23 83 24
rect 83 23 84 24
rect 84 23 85 24
rect 85 23 86 24
rect 86 23 87 24
rect 87 23 88 24
rect 88 23 89 24
rect 89 23 90 24
rect 90 23 91 24
rect 91 23 92 24
rect 92 23 93 24
rect 93 23 94 24
rect 94 23 95 24
rect 95 23 96 24
rect 96 23 97 24
rect 97 23 98 24
rect 98 23 99 24
rect 99 23 100 24
rect 100 23 101 24
rect 101 23 102 24
rect 102 23 103 24
rect 103 23 104 24
rect 104 23 105 24
rect 105 23 106 24
rect 106 23 107 24
rect 107 23 108 24
rect 108 23 109 24
rect 109 23 110 24
rect 110 23 111 24
rect 111 23 112 24
rect 112 23 113 24
rect 113 23 114 24
rect 114 23 115 24
rect 115 23 116 24
rect 116 23 117 24
rect 117 23 118 24
rect 118 23 119 24
rect 119 23 120 24
rect 120 23 121 24
rect 121 23 122 24
rect 122 23 123 24
rect 123 23 124 24
rect 124 23 125 24
rect 125 23 126 24
rect 126 23 127 24
rect 127 23 128 24
rect 128 23 129 24
rect 129 23 130 24
rect 130 23 131 24
rect 131 23 132 24
rect 132 23 133 24
rect 133 23 134 24
rect 134 23 135 24
rect 164 23 165 24
rect 165 23 166 24
rect 166 23 167 24
rect 167 23 168 24
rect 168 23 169 24
rect 169 23 170 24
rect 83 22 84 23
rect 84 22 85 23
rect 85 22 86 23
rect 86 22 87 23
rect 87 22 88 23
rect 88 22 89 23
rect 89 22 90 23
rect 90 22 91 23
rect 91 22 92 23
rect 92 22 93 23
rect 93 22 94 23
rect 94 22 95 23
rect 95 22 96 23
rect 96 22 97 23
rect 97 22 98 23
rect 98 22 99 23
rect 99 22 100 23
rect 100 22 101 23
rect 101 22 102 23
rect 102 22 103 23
rect 103 22 104 23
rect 104 22 105 23
rect 105 22 106 23
rect 106 22 107 23
rect 107 22 108 23
rect 108 22 109 23
rect 109 22 110 23
rect 110 22 111 23
rect 111 22 112 23
rect 112 22 113 23
rect 113 22 114 23
rect 114 22 115 23
rect 115 22 116 23
rect 116 22 117 23
rect 117 22 118 23
rect 118 22 119 23
rect 119 22 120 23
rect 120 22 121 23
rect 121 22 122 23
rect 122 22 123 23
rect 123 22 124 23
rect 124 22 125 23
rect 125 22 126 23
rect 126 22 127 23
rect 127 22 128 23
rect 128 22 129 23
rect 129 22 130 23
rect 130 22 131 23
rect 131 22 132 23
rect 132 22 133 23
rect 133 22 134 23
rect 163 22 164 23
rect 164 22 165 23
rect 165 22 166 23
rect 166 22 167 23
rect 167 22 168 23
rect 168 22 169 23
rect 85 21 86 22
rect 86 21 87 22
rect 87 21 88 22
rect 88 21 89 22
rect 89 21 90 22
rect 90 21 91 22
rect 91 21 92 22
rect 92 21 93 22
rect 93 21 94 22
rect 94 21 95 22
rect 95 21 96 22
rect 96 21 97 22
rect 97 21 98 22
rect 98 21 99 22
rect 99 21 100 22
rect 100 21 101 22
rect 101 21 102 22
rect 102 21 103 22
rect 103 21 104 22
rect 104 21 105 22
rect 105 21 106 22
rect 106 21 107 22
rect 107 21 108 22
rect 108 21 109 22
rect 109 21 110 22
rect 110 21 111 22
rect 111 21 112 22
rect 112 21 113 22
rect 113 21 114 22
rect 114 21 115 22
rect 115 21 116 22
rect 116 21 117 22
rect 117 21 118 22
rect 118 21 119 22
rect 119 21 120 22
rect 120 21 121 22
rect 121 21 122 22
rect 122 21 123 22
rect 123 21 124 22
rect 124 21 125 22
rect 125 21 126 22
rect 126 21 127 22
rect 127 21 128 22
rect 128 21 129 22
rect 129 21 130 22
rect 130 21 131 22
rect 131 21 132 22
rect 132 21 133 22
rect 133 21 134 22
rect 161 21 162 22
rect 162 21 163 22
rect 163 21 164 22
rect 164 21 165 22
rect 165 21 166 22
rect 166 21 167 22
rect 167 21 168 22
rect 87 20 88 21
rect 88 20 89 21
rect 89 20 90 21
rect 90 20 91 21
rect 91 20 92 21
rect 92 20 93 21
rect 93 20 94 21
rect 94 20 95 21
rect 95 20 96 21
rect 96 20 97 21
rect 97 20 98 21
rect 98 20 99 21
rect 99 20 100 21
rect 100 20 101 21
rect 101 20 102 21
rect 102 20 103 21
rect 103 20 104 21
rect 104 20 105 21
rect 105 20 106 21
rect 106 20 107 21
rect 107 20 108 21
rect 108 20 109 21
rect 109 20 110 21
rect 110 20 111 21
rect 111 20 112 21
rect 112 20 113 21
rect 113 20 114 21
rect 114 20 115 21
rect 115 20 116 21
rect 116 20 117 21
rect 117 20 118 21
rect 118 20 119 21
rect 119 20 120 21
rect 120 20 121 21
rect 121 20 122 21
rect 122 20 123 21
rect 123 20 124 21
rect 124 20 125 21
rect 125 20 126 21
rect 126 20 127 21
rect 127 20 128 21
rect 128 20 129 21
rect 129 20 130 21
rect 130 20 131 21
rect 131 20 132 21
rect 132 20 133 21
rect 133 20 134 21
rect 134 20 135 21
rect 135 20 136 21
rect 160 20 161 21
rect 161 20 162 21
rect 162 20 163 21
rect 163 20 164 21
rect 164 20 165 21
rect 165 20 166 21
rect 166 20 167 21
rect 88 19 89 20
rect 89 19 90 20
rect 90 19 91 20
rect 91 19 92 20
rect 92 19 93 20
rect 93 19 94 20
rect 94 19 95 20
rect 95 19 96 20
rect 96 19 97 20
rect 97 19 98 20
rect 98 19 99 20
rect 99 19 100 20
rect 100 19 101 20
rect 101 19 102 20
rect 102 19 103 20
rect 103 19 104 20
rect 104 19 105 20
rect 105 19 106 20
rect 106 19 107 20
rect 107 19 108 20
rect 108 19 109 20
rect 109 19 110 20
rect 110 19 111 20
rect 111 19 112 20
rect 112 19 113 20
rect 113 19 114 20
rect 114 19 115 20
rect 115 19 116 20
rect 116 19 117 20
rect 117 19 118 20
rect 118 19 119 20
rect 119 19 120 20
rect 120 19 121 20
rect 121 19 122 20
rect 122 19 123 20
rect 123 19 124 20
rect 124 19 125 20
rect 125 19 126 20
rect 126 19 127 20
rect 127 19 128 20
rect 128 19 129 20
rect 129 19 130 20
rect 130 19 131 20
rect 131 19 132 20
rect 132 19 133 20
rect 133 19 134 20
rect 134 19 135 20
rect 135 19 136 20
rect 136 19 137 20
rect 158 19 159 20
rect 159 19 160 20
rect 160 19 161 20
rect 161 19 162 20
rect 162 19 163 20
rect 163 19 164 20
rect 164 19 165 20
rect 90 18 91 19
rect 91 18 92 19
rect 92 18 93 19
rect 93 18 94 19
rect 94 18 95 19
rect 95 18 96 19
rect 96 18 97 19
rect 97 18 98 19
rect 98 18 99 19
rect 99 18 100 19
rect 100 18 101 19
rect 101 18 102 19
rect 102 18 103 19
rect 103 18 104 19
rect 104 18 105 19
rect 105 18 106 19
rect 106 18 107 19
rect 107 18 108 19
rect 108 18 109 19
rect 109 18 110 19
rect 110 18 111 19
rect 111 18 112 19
rect 112 18 113 19
rect 113 18 114 19
rect 114 18 115 19
rect 115 18 116 19
rect 116 18 117 19
rect 117 18 118 19
rect 118 18 119 19
rect 119 18 120 19
rect 120 18 121 19
rect 121 18 122 19
rect 122 18 123 19
rect 123 18 124 19
rect 124 18 125 19
rect 125 18 126 19
rect 126 18 127 19
rect 127 18 128 19
rect 128 18 129 19
rect 129 18 130 19
rect 130 18 131 19
rect 131 18 132 19
rect 132 18 133 19
rect 133 18 134 19
rect 134 18 135 19
rect 135 18 136 19
rect 136 18 137 19
rect 137 18 138 19
rect 138 18 139 19
rect 139 18 140 19
rect 140 18 141 19
rect 153 18 154 19
rect 154 18 155 19
rect 155 18 156 19
rect 156 18 157 19
rect 157 18 158 19
rect 158 18 159 19
rect 159 18 160 19
rect 160 18 161 19
rect 161 18 162 19
rect 162 18 163 19
rect 163 18 164 19
rect 164 18 165 19
rect 112 17 113 18
rect 113 17 114 18
rect 114 17 115 18
rect 115 17 116 18
rect 116 17 117 18
rect 117 17 118 18
rect 118 17 119 18
rect 119 17 120 18
rect 120 17 121 18
rect 121 17 122 18
rect 122 17 123 18
rect 123 17 124 18
rect 124 17 125 18
rect 125 17 126 18
rect 126 17 127 18
rect 127 17 128 18
rect 128 17 129 18
rect 129 17 130 18
rect 130 17 131 18
rect 131 17 132 18
rect 132 17 133 18
rect 133 17 134 18
rect 134 17 135 18
rect 135 17 136 18
rect 136 17 137 18
rect 137 17 138 18
rect 138 17 139 18
rect 139 17 140 18
rect 140 17 141 18
rect 141 17 142 18
rect 142 17 143 18
rect 143 17 144 18
rect 144 17 145 18
rect 145 17 146 18
rect 146 17 147 18
rect 149 17 150 18
rect 150 17 151 18
rect 151 17 152 18
rect 152 17 153 18
rect 153 17 154 18
rect 154 17 155 18
rect 155 17 156 18
rect 156 17 157 18
rect 157 17 158 18
rect 158 17 159 18
rect 159 17 160 18
rect 160 17 161 18
rect 161 17 162 18
rect 115 16 116 17
rect 116 16 117 17
rect 117 16 118 17
rect 118 16 119 17
rect 119 16 120 17
rect 120 16 121 17
rect 121 16 122 17
rect 122 16 123 17
rect 123 16 124 17
rect 124 16 125 17
rect 125 16 126 17
rect 126 16 127 17
rect 127 16 128 17
rect 128 16 129 17
rect 129 16 130 17
rect 130 16 131 17
rect 131 16 132 17
rect 132 16 133 17
rect 133 16 134 17
rect 134 16 135 17
rect 135 16 136 17
rect 136 16 137 17
rect 137 16 138 17
rect 138 16 139 17
rect 139 16 140 17
rect 140 16 141 17
rect 141 16 142 17
rect 142 16 143 17
rect 143 16 144 17
rect 144 16 145 17
rect 145 16 146 17
rect 146 16 147 17
rect 147 16 148 17
rect 148 16 149 17
rect 149 16 150 17
rect 150 16 151 17
rect 151 16 152 17
rect 152 16 153 17
rect 153 16 154 17
rect 154 16 155 17
rect 155 16 156 17
rect 156 16 157 17
rect 157 16 158 17
rect 158 16 159 17
rect 159 16 160 17
rect 160 16 161 17
rect 118 15 119 16
rect 119 15 120 16
rect 120 15 121 16
rect 121 15 122 16
rect 122 15 123 16
rect 123 15 124 16
rect 124 15 125 16
rect 125 15 126 16
rect 126 15 127 16
rect 127 15 128 16
rect 128 15 129 16
rect 129 15 130 16
rect 130 15 131 16
rect 131 15 132 16
rect 132 15 133 16
rect 133 15 134 16
rect 134 15 135 16
rect 135 15 136 16
rect 136 15 137 16
rect 137 15 138 16
rect 138 15 139 16
rect 139 15 140 16
rect 140 15 141 16
rect 141 15 142 16
rect 142 15 143 16
rect 143 15 144 16
rect 144 15 145 16
rect 145 15 146 16
rect 146 15 147 16
rect 147 15 148 16
rect 148 15 149 16
rect 149 15 150 16
rect 150 15 151 16
rect 151 15 152 16
rect 152 15 153 16
rect 153 15 154 16
rect 154 15 155 16
rect 155 15 156 16
rect 156 15 157 16
rect 157 15 158 16
rect 158 15 159 16
rect 159 15 160 16
rect 120 14 121 15
rect 121 14 122 15
rect 122 14 123 15
rect 123 14 124 15
rect 124 14 125 15
rect 125 14 126 15
rect 126 14 127 15
rect 127 14 128 15
rect 128 14 129 15
rect 129 14 130 15
rect 130 14 131 15
rect 131 14 132 15
rect 132 14 133 15
rect 133 14 134 15
rect 134 14 135 15
rect 135 14 136 15
rect 136 14 137 15
rect 137 14 138 15
rect 138 14 139 15
rect 139 14 140 15
rect 140 14 141 15
rect 141 14 142 15
rect 142 14 143 15
rect 143 14 144 15
rect 144 14 145 15
rect 145 14 146 15
rect 146 14 147 15
rect 147 14 148 15
rect 148 14 149 15
rect 149 14 150 15
rect 150 14 151 15
rect 151 14 152 15
rect 152 14 153 15
rect 153 14 154 15
rect 154 14 155 15
rect 155 14 156 15
rect 156 14 157 15
rect 157 14 158 15
rect 158 14 159 15
rect 123 13 124 14
rect 124 13 125 14
rect 125 13 126 14
rect 126 13 127 14
rect 127 13 128 14
rect 128 13 129 14
rect 129 13 130 14
rect 130 13 131 14
rect 131 13 132 14
rect 132 13 133 14
rect 133 13 134 14
rect 134 13 135 14
rect 135 13 136 14
rect 136 13 137 14
rect 137 13 138 14
rect 138 13 139 14
rect 139 13 140 14
rect 140 13 141 14
rect 141 13 142 14
rect 142 13 143 14
rect 143 13 144 14
rect 144 13 145 14
rect 145 13 146 14
rect 146 13 147 14
rect 147 13 148 14
rect 148 13 149 14
rect 149 13 150 14
rect 150 13 151 14
rect 151 13 152 14
rect 152 13 153 14
rect 153 13 154 14
rect 154 13 155 14
rect 155 13 156 14
rect 156 13 157 14
rect 125 12 126 13
rect 126 12 127 13
rect 127 12 128 13
rect 128 12 129 13
rect 129 12 130 13
rect 130 12 131 13
rect 131 12 132 13
rect 132 12 133 13
rect 133 12 134 13
rect 134 12 135 13
rect 135 12 136 13
rect 136 12 137 13
rect 137 12 138 13
rect 138 12 139 13
rect 139 12 140 13
rect 140 12 141 13
rect 141 12 142 13
rect 142 12 143 13
rect 143 12 144 13
rect 144 12 145 13
rect 145 12 146 13
rect 146 12 147 13
rect 147 12 148 13
rect 148 12 149 13
rect 149 12 150 13
rect 150 12 151 13
rect 151 12 152 13
rect 152 12 153 13
rect 153 12 154 13
rect 154 12 155 13
rect 155 12 156 13
rect 156 12 157 13
rect 128 11 129 12
rect 129 11 130 12
rect 130 11 131 12
rect 131 11 132 12
rect 132 11 133 12
rect 133 11 134 12
rect 134 11 135 12
rect 135 11 136 12
rect 136 11 137 12
rect 137 11 138 12
rect 138 11 139 12
rect 139 11 140 12
rect 140 11 141 12
rect 141 11 142 12
rect 142 11 143 12
rect 143 11 144 12
rect 144 11 145 12
rect 145 11 146 12
rect 146 11 147 12
rect 147 11 148 12
rect 148 11 149 12
rect 149 11 150 12
rect 150 11 151 12
rect 151 11 152 12
rect 152 11 153 12
rect 153 11 154 12
rect 154 11 155 12
rect 132 10 133 11
rect 133 10 134 11
rect 134 10 135 11
rect 135 10 136 11
rect 136 10 137 11
rect 137 10 138 11
rect 138 10 139 11
rect 139 10 140 11
rect 140 10 141 11
rect 141 10 142 11
rect 142 10 143 11
rect 143 10 144 11
rect 144 10 145 11
rect 145 10 146 11
rect 146 10 147 11
rect 147 10 148 11
rect 148 10 149 11
rect 149 10 150 11
rect 150 10 151 11
rect 151 10 152 11
rect 152 10 153 11
rect 136 9 137 10
rect 137 9 138 10
rect 138 9 139 10
rect 139 9 140 10
rect 140 9 141 10
rect 141 9 142 10
rect 142 9 143 10
rect 143 9 144 10
rect 144 9 145 10
rect 145 9 146 10
rect 146 9 147 10
rect 147 9 148 10
rect 148 9 149 10
rect 149 9 150 10
rect 150 9 151 10
rect 151 9 152 10
rect 140 8 141 9
rect 141 8 142 9
rect 142 8 143 9
rect 143 8 144 9
rect 144 8 145 9
rect 145 8 146 9
rect 146 8 147 9
rect 147 8 148 9
rect 148 8 149 9
rect 149 8 150 9
rect 150 8 151 9
<< end >>
