VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO comp_a
  CLASS BLOCK ;
  FOREIGN comp_a ;
  ORIGIN 0.000 0.000 ;
  SIZE 10000.000 BY 2000.000 ;
END comp_a
END LIBRARY

