* Extracted by KLayout

* cell testall
.SUBCKT testall
* cell instance $2 r0 *1 0,0
X$2 1 2 FDPTEST
* cell instance $3 r0 *1 0,0
X$3 4 1 FWBTEST
* cell instance $7 r0 *1 0,0
X$7 5 1 DPTEST
* cell instance $8 r0 *1 0,0
X$8 2 3 FBGATEST
* cell instance $9 r0 *1 0,0
X$9 5 6 BDPTEST
* cell instance $10 r0 *1 0,0
X$10 8 5 BWBTEST
* cell instance $14 r0 *1 0,0
X$14 7 6 BBGATEST
.ENDS testall

* cell FDPTEST
* pin B
* pin A
.SUBCKT FDPTEST 1 2
.ENDS FDPTEST

* cell DPTEST
* pin B
* pin A
.SUBCKT DPTEST 1 2
.ENDS DPTEST

* cell BDPTEST
* pin A
* pin B
.SUBCKT BDPTEST 1 2
.ENDS BDPTEST

* cell BBGATEST
* pin B
* pin A
.SUBCKT BBGATEST 1 2
.ENDS BBGATEST

* cell FBGATEST
* pin B
* pin A
.SUBCKT FBGATEST 1 2
.ENDS FBGATEST

* cell FWBTEST
* pin B
* pin A
.SUBCKT FWBTEST 1 2
.ENDS FWBTEST

* cell BWBTEST
* pin B
* pin A
.SUBCKT BWBTEST 1 2
.ENDS BWBTEST
