* Extracted by KLayout

.SUBCKT TOP A Q VDD SUBSTRATE|VSS
X$1 SUBSTRATE|VSS VDD VDD \$1 Q SUBSTRATE|VSS INV
X$2 SUBSTRATE|VSS VDD VDD A \$1 SUBSTRATE|VSS INV
.ENDS TOP

.SUBCKT INV \$1 \$2 \$3 \$4 \$5 SUBSTRATE
X$1 \$5 \$1 \$4 SUBSTRATE NTRANS
X$2 \$5 \$2 \$4 \$3 PTRANS
.ENDS INV

.SUBCKT NTRANS \$1 \$3 \$5 SUBSTRATE
M$1 \$3 \$5 \$1 SUBSTRATE NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
.ENDS NTRANS

.SUBCKT PTRANS \$1 \$3 \$5 \$I3
M$1 \$3 \$5 \$1 \$I3 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
.ENDS PTRANS
