* Extracted by KLayout

* cell testall
.SUBCKT testall
* cell instance $2 r0 *1 0,0
X$2 1 3 FDPTEST
* cell instance $3 r0 *1 0,0
X$3 1 FWBTEST
* cell instance $7 r0 *1 0,0
X$7 2 1 DPTEST
* cell instance $8 r0 *1 0,0
X$8 2 2 BDPTEST
* cell instance $9 r0 *1 0,0
X$9 2 BBGATEST
* cell instance $10 r0 *1 0,0
X$10 2 BWBTEST
* cell instance $14 r0 *1 0,0
X$14 3 FBGATEST
.ENDS testall

* cell FDPTEST
* pin B
* pin A
.SUBCKT FDPTEST 1 2
* net 1 B
* net 2 A
.ENDS FDPTEST

* cell DPTEST
* pin B
* pin A
.SUBCKT DPTEST 1 2
* net 1 B
* net 2 A
.ENDS DPTEST

* cell BDPTEST
* pin A
* pin B
.SUBCKT BDPTEST 1 2
* net 1 A
* net 2 B
.ENDS BDPTEST

* cell BBGATEST
* pin A
.SUBCKT BBGATEST 2
* net 1 B
* net 2 A
.ENDS BBGATEST

* cell FBGATEST
* pin B
.SUBCKT FBGATEST 1
* net 1 B
* net 2 A
.ENDS FBGATEST

* cell FWBTEST
* pin A
.SUBCKT FWBTEST 2
* net 1 B
* net 2 A
.ENDS FWBTEST

* cell BWBTEST
* pin A
.SUBCKT BWBTEST 2
* net 1 B
* net 2 A
.ENDS BWBTEST
