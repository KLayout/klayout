magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 540 108 756
rect 0 504 252 540
rect 0 468 288 504
rect 0 396 324 468
rect 0 0 108 396
rect 216 0 324 396
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
