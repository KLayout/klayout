magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 6300 6120 6804 6156
rect 6264 6084 6840 6120
rect 6228 6048 6876 6084
rect 6192 6012 6372 6048
rect 6732 6012 6912 6048
rect 6156 5976 6336 6012
rect 6768 5976 6912 6012
rect 6156 5940 6300 5976
rect 6156 5400 6264 5940
rect 6444 5904 6624 5940
rect 6408 5868 6660 5904
rect 6372 5796 6696 5868
rect 6372 5544 6480 5796
rect 6588 5724 6696 5796
rect 6588 5544 6696 5616
rect 6372 5472 6696 5544
rect 6408 5436 6660 5472
rect 6444 5400 6624 5436
rect 6804 5400 6912 5976
rect 6156 5364 6300 5400
rect 6768 5364 6912 5400
rect 6156 5328 6336 5364
rect 6732 5328 6912 5364
rect 6192 5292 6372 5328
rect 6696 5292 6876 5328
rect 6228 5256 6840 5292
rect 6264 5220 6804 5256
rect 6300 5184 6768 5220
<< end >>
