
VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
USEMINSPACING OBS OFF ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  OFFSET 0.17 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;
  SPACING 0.17 ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  OFFSET 0.23 ;
  WIDTH 0.14 ; 
END met2

LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ; 
  SPACING 0.2 ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  OFFSET 0.34 ;
  WIDTH 0.3 ; 
END met3

VIA via1 DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.24 0.16 0.24 ;
  LAYER met2 ;
  RECT -0.13 -0.24 0.13 0.24 ;
END via1

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

VIA via2 DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.24 0.14 0.24 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END via2

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

END LIBRARY
 
