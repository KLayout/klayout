
* Simple CMOS inverer circuit 

.SUBCKT INVERTER_WITH_DIODES VSS IN OUT VDD 
Mp VDD IN OUT VDD PMOS W=1.5U L=0.25U
Mn OUT IN VSS VSS NMOS W=0.9U L=0.25U
.ENDS

