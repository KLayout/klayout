
* cell LVS_TEST
* pin VDDO
* pin VP
.SUBCKT LVS_TEST 1 2
* net 1 VDDO
* net 2 VP
* device instance 1I38 r0 *1 0,0 PCH_18_MAC
M1I38 1 2 1 1 PCH_18_MAC L=0.225U W=10653U AS=0P AD=0P PS=0U PD=0U
* device instance 1I39A r0 *1 0,0 PCH_18_MAC
M1I39A 1 2 1 1 PCH_18_MAC L=0.135U W=1809U AS=0P AD=0P PS=0U PD=0U
.ENDS LVS_TEST
