
.SUBCKT XPMOS S G D B PARAMS: L=1U W=1U
  M$1 S G D B PMOS L=L W=W
.ENDS PMOS

.SUBCKT NMOS S G D B PARAMS: L=1U W=1U
  M$1 S G D B NMOS L=L W=W
.ENDS NMOS

.SUBCKT RINGO VSS VDD FB ENABLE OUT
X$1 VDD 1 VSS VDD FB ENABLE VSS ND2X1
X$2 VDD 2 VSS VDD 1 VSS INVX1
X$3 VDD 3 VSS VDD 2 VSS INVX1
X$4 VDD 4 VSS VDD 3 VSS INVX1
X$5 VDD 5 VSS VDD 4 VSS INVX1
X$6 VDD 6 VSS VDD 5 VSS INVX1
X$7 VDD 7 VSS VDD 6 VSS INVX1
X$8 VDD 8 VSS VDD 7 VSS INVX1
X$9 VDD 9 VSS VDD 8 VSS INVX1
X$10 VDD 10 VSS VDD 9 VSS INVX1
X$11 VDD FB VSS VDD 10 VSS INVX1
X$12 VDD OUT VSS VDD FB VSS INVX1
.ENDS RINGO

.SUBCKT ND2X1 VDD OUT VSS NWELL B A BULK
X$1 OUT A VDD NWELL XPMOS L=0.25U W=1.5U 
X$2 VDD B OUT NWELL XPMOS L=0.25U W=1.5U 
X$3 VSS A 1 BULK NMOS L=0.25U W=0.95U 
X$4 1 B OUT BULK NMOS L=0.25U W=0.95U 
.ENDS ND2X1

.SUBCKT INVX1 VDD OUT VSS NWELL IN BULK
X$1 VDD IN OUT NWELL XPMOS L=0.25U W=1.5U 
X$2 VSS IN OUT BULK NMOS L=0.25U W=0.95U 
.ENDS INVX1
