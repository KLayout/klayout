* RINGO netlist before simplification

* cell RINGO
.SUBCKT RINGO
* net 12 OUT
* net 27 ENABLE
* net 28 VDD
* net 29 FB
* net 43 BULK,VSS
* device instance $1 2.65,5.8 LVPMOS
M$1 2 27 28 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 3.35,5.8 LVPMOS
M$2 28 29 2 28 LVPMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 5.05,5.8 LVPMOS
M$3 28 2 3 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $4 6.85,5.8 LVPMOS
M$4 28 3 4 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $5 8.65,5.8 LVPMOS
M$5 28 4 5 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $6 10.45,5.8 LVPMOS
M$6 28 5 6 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $7 12.25,5.8 LVPMOS
M$7 28 6 7 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $8 14.05,5.8 LVPMOS
M$8 28 7 8 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $9 15.85,5.8 LVPMOS
M$9 28 8 9 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $10 17.65,5.8 LVPMOS
M$10 28 9 10 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $11 19.45,5.8 LVPMOS
M$11 28 10 11 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $12 21.25,5.8 LVPMOS
M$12 28 11 29 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $13 23.05,5.8 LVPMOS
M$13 28 29 12 28 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $14 2.65,2.135 LVNMOS
M$14 43 27 14 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U
+ PD=1.4U
* device instance $15 3.35,2.135 LVNMOS
M$15 14 29 2 43 LVNMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
* device instance $16 5.05,2.135 LVNMOS
M$16 43 2 3 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $17 6.85,2.135 LVNMOS
M$17 43 3 4 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $18 8.65,2.135 LVNMOS
M$18 43 4 5 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $19 10.45,2.135 LVNMOS
M$19 43 5 6 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $20 12.25,2.135 LVNMOS
M$20 43 6 7 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $21 14.05,2.135 LVNMOS
M$21 43 7 8 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $22 15.85,2.135 LVNMOS
M$22 43 8 9 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $23 17.65,2.135 LVNMOS
M$23 43 9 10 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
* device instance $24 19.45,2.135 LVNMOS
M$24 43 10 11 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
* device instance $25 21.25,2.135 LVNMOS
M$25 43 11 29 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
* device instance $26 23.05,2.135 LVNMOS
M$26 43 29 12 43 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
.ENDS RINGO
