* VDIV netlist before simplification

* cell TOP
.SUBCKT TOP
* net 1 OUT
* net 2 GND
* net 4 IN
* net 7 VDD
* device instance $1 1.025,0.335 RES
R$1 6 1 7650
* device instance $2 2.85,0.335 RES
R$2 3 1 7650
* device instance $3 4.665,0.335 RES
R$3 3 2 2670
* device instance $4 1.765,7.485 HVPMOS
M$4 6 4 7 7 HVPMOS L=0.25U W=1.5U AS=0.63P AD=0.63P PS=3.84U PD=3.84U
.ENDS TOP
