magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 720 144 756
rect 0 684 180 720
rect 0 612 216 684
rect 108 504 216 612
rect 108 432 252 504
rect 144 324 324 432
rect 108 252 252 324
rect 108 144 216 252
rect 0 72 216 144
rect 0 36 180 72
rect 0 0 144 36
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
