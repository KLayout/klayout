magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 648 108 756
rect 0 540 216 648
rect 324 540 432 756
rect 0 432 432 540
rect 0 0 108 432
rect 216 324 432 432
rect 324 0 432 324
<< properties >>
string FIXED_BBOX 0 -216 540 756
<< end >>
