VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
  LAYER LEF58_MINWIDTH STRING ; 
END PROPERTYDEFINITIONS

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
    WIDTH 0.6 ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
    WIDTH 0.5 ;
       PROPERTY LEF58_MINWIDTH "MINWIDTH 1.0 WRONGDIRECTION ; " ;
END M4

VIA via34
	LAYER M3 ; 
		RECT -0.4 -0.3 0.4 0.3 ;
	LAYER VIA3 ; 
		RECT -0.3 -0.25 0.3 0.25 ;
	LAYER M4 ;
		RECT -1.00 -0.5 1.00 0.5 ;
END via34

END LIBRARY
