.SUBCKT INV_CHAIN 1 2
M2_1.N1 4 3 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_1.P1 4 3 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_2.N1 5 4 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_2.P1 5 4 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_3.N1 6 5 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_3.P1 6 5 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_4.N1 7 6 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_4.P1 7 6 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_5.N1 8 7 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M2_5.P1 8 7 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_1.N1 10 9 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_1.P1 10 9 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_2.N1 11 10 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_2.P1 11 10 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_3.N1 12 11 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_3.P1 12 11 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_4.N1 13 12 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_4.P1 13 12 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_5.N1 14 13 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M_5.P1 14 13 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_1.N1 16 15 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_1.P1 16 15 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_2.N1 17 16 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_2.P1 17 16 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_3.N1 18 17 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_3.P1 18 17 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_4.N1 19 18 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_4.P1 19 18 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_5.N1 20 19 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_5.P1 20 19 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_6.N1 21 20 2 2 NCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
M0_6.P1 21 20 1 1 PCH_SVT_MAC L=0.016U W=3U AS=0P AD=0P PS=0U PD=0U
.ENDS INV_CHAIN
