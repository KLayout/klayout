magic
tech scmos
timestamp 1534225390
<< silk >>
rect 0 4 4 18
rect 8 4 12 6
rect 0 0 12 4
<< end >>
