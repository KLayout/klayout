* RINGO netlist with global nets

.GLOBAL VDD
.GLOBAL VSS

.SUBCKT RINGO FB OUT ENABLE 
X$1 1 FB ENABLE ND2X1
X$2 2 1 INVX1
X$3 3 2 INVX1
X$4 4 3 INVX1
X$5 5 4 INVX1
X$6 6 5 INVX1
X$7 7 6 INVX1
X$8 8 7 INVX1
X$9 9 8 INVX1
X$10 10 9 INVX1
X$11 FB 10 INVX1
X$12 OUT FB INVX1
.ENDS RINGO

.SUBCKT ND2X1 OUT B A 
M$1 OUT A VDD VDD MLVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
M$2 VDD B OUT VDD MLVPMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
M$3 VSS A INT VSS MLVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U PD=1.4U
M$4 INT B OUT VSS MLVNMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
.ENDS ND2X1

.SUBCKT INVX1 OUT IN 
M$1 VDD IN OUT VDD MLVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
M$2 VSS IN OUT VSS MLVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
.ENDS INVX1
