magic
tech scmos
timestamp 1534325697
<< silk >>
rect 0 0 4 4
<< end >>
