magic
tech scmos
timestamp 1534322005
<< silk >>
rect 2 17 10 18
rect 1 16 11 17
rect 0 14 12 16
rect 0 4 4 14
rect 8 13 12 14
rect 7 7 12 10
rect 9 4 12 7
rect 0 3 5 4
rect 8 3 12 4
rect 0 2 12 3
rect 1 1 12 2
rect 2 0 12 1
<< end >>
