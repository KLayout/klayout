magic
tech scmos
timestamp 1533654616
<< pwell >>
rect 0 0 24 23
<< nwell >>
rect 0 32 24 56
<< polysilicon >>
rect 7 46 9 48
rect 15 46 17 48
rect 7 33 9 35
rect 15 33 17 35
rect 7 32 17 33
rect 7 31 10 32
rect 14 31 17 32
rect 6 24 9 25
rect 3 23 9 24
rect 7 21 9 23
rect 15 24 18 25
rect 15 23 21 24
rect 15 21 17 23
rect 7 8 9 10
rect 15 8 17 10
<< ndiffusion >>
rect 6 10 7 21
rect 9 10 10 21
rect 14 10 15 21
rect 17 10 18 21
<< pdiffusion >>
rect 6 35 7 46
rect 9 35 10 46
rect 14 35 15 46
rect 17 35 18 46
<< metal1 >>
rect 0 50 2 54
rect 22 50 24 54
rect 10 46 14 50
rect 2 28 6 35
rect 10 21 14 28
rect 18 28 22 35
rect 2 6 6 10
rect 18 6 22 10
rect 0 2 2 6
rect 22 2 24 6
<< ntransistor >>
rect 7 10 9 21
rect 15 10 17 21
<< ptransistor >>
rect 7 35 9 46
rect 15 35 17 46
<< polycontact >>
rect 10 28 14 32
rect 2 24 6 28
rect 18 24 22 28
<< ndcontact >>
rect 2 10 6 21
rect 10 10 14 21
rect 18 10 22 21
<< pdcontact >>
rect 2 35 6 46
rect 10 35 14 46
rect 18 35 22 46
<< psubstratepcontact >>
rect 2 2 22 6
<< nsubstratencontact >>
rect 2 50 22 54
<< labels >>
rlabel psubstratepcontact 2 2 22 6 1 gnd!
rlabel nsubstratencontact 2 50 22 54 1 vdd!
<< end >>
