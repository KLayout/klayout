* Extracted by KLayout

* cell RINGO
* pin FB
* pin VDD
* pin OUT
* pin ENABLE
* pin VSS
.SUBCKT RINGO 12 13 14 15 16
* net 12 FB
* net 13 VDD
* net 14 OUT
* net 15 ENABLE
* net 16 VSS
* cell instance $3 r0 *1 1.8,0
X$3 13 2 16 13 12 15 16 ND2X1
* cell instance $4 r0 *1 4.2,0
X$4 13 3 16 13 2 16 INVX1
* cell instance $5 r0 *1 6,0
X$5 13 4 16 13 3 16 INVX1
* cell instance $6 r0 *1 7.8,0
X$6 13 5 16 13 4 16 INVX1
* cell instance $7 r0 *1 9.6,0
X$7 13 6 16 13 5 16 INVX1
* cell instance $8 r0 *1 11.4,0
X$8 13 7 16 13 6 16 INVX1
* cell instance $9 r0 *1 13.2,0
X$9 13 8 16 13 7 16 INVX1
* cell instance $10 r0 *1 15,0
X$10 13 9 16 13 8 16 INVX1
* cell instance $11 r0 *1 16.8,0
X$11 13 10 16 13 9 16 INVX1
* cell instance $12 r0 *1 18.6,0
X$12 13 11 16 13 10 16 INVX1
* cell instance $13 r0 *1 20.4,0
X$13 13 12 16 13 11 16 INVX1
* cell instance $14 r0 *1 22.2,0
X$14 13 14 16 13 12 16 INVX1
* device instance $1 r0 *1 26.45,2.075 NMOS
M$1 16 1 16 16 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
.ENDS RINGO

* cell INVX1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin IN
* pin SUBSTRATE
.SUBCKT INVX1 1 2 3 4 5 6
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 IN
* net 6 SUBSTRATE
* device instance $1 r0 *1 0.85,5.8 PMOS
M$1 1 5 2 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $2 r0 *1 0.85,2.135 NMOS
M$2 3 5 2 6 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
.ENDS INVX1

* cell ND2X1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin B
* pin A
* pin SUBSTRATE
.SUBCKT ND2X1 1 2 3 4 5 6 7
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 B
* net 6 A
* net 7 SUBSTRATE
* device instance $1 r0 *1 0.85,5.8 PMOS
M$1 2 6 1 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 r0 *1 1.55,5.8 PMOS
M$2 1 5 2 4 PMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 r0 *1 0.85,2.135 NMOS
M$3 3 6 8 7 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U PD=1.4U
* device instance $4 r0 *1 1.55,2.135 NMOS
M$4 8 5 2 7 NMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
.ENDS ND2X1
