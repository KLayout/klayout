VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

LAYER mx
    TYPE ROUTING ;
    WIDTH 0.04 ;
    DIRECTION HORIZONTAL ;
    PROPERTY LEF58_WIDTHTABLE "
      WIDTHTABLE 0.08  ;
      WIDTHTABLE 0.12 WRONGDIRECTION ;
    " ;
END mx
END LIBRARY
