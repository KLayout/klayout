VERSION 5.8 ;

MACRO a
  ORIGIN 0 0 ;
  SIZE 600 BY 600 ;
  OBS 
    LAYER M1 ;
      RECT 10 10 590 590 ;
  END
END a

MACRO b
  ORIGIN -600 0 ;
  SIZE 400 BY 500 ;
  OBS 
    LAYER M1 ;
      RECT 610 10 990 490 ;
  END
END b

MACRO c
  ORIGIN -500 -500 ;
  SIZE 500 BY 500 ;
  OBS 
    LAYER M1 ;
      POLYGON 510 610 610 610 610 510 990 510 990 990 510 990 ;
    LAYER overlap ;
      RECT 500 700 1000 1000 ;
      POLYGON 500 600  600 600  600 500  1000 500  1000 700  500 700 ;
  END
END c
