magic
tech scmos
timestamp 1534321628
<< silk >>
rect 0 16 10 18
rect 0 14 12 16
rect 0 11 4 14
rect 7 11 12 14
rect 0 8 11 11
rect 0 4 4 8
rect 8 5 12 8
rect 7 4 12 5
rect 0 2 12 4
rect 0 0 10 2
<< end >>
