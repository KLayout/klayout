
.SUBCKT RINGO VSS VDD FB ENABLE OUT
X$1 VDD VSS 1 FB ENABLE ND2X1
X$2 VDD VSS 2 1 INVX1
X$3 VDD VSS 3 2 INVX1
X$4 VDD VSS 4 3 INVX1
X$5 VDD VSS 5 4 INVX1
X$6 VDD VSS 6 5 INVX1
X$7 VDD VSS 7 6 INVX1
X$8 VDD VSS 8 7 INVX1
X$9 VDD VSS 9 8 INVX1
X$10 VDD VSS 10 9 INVX1
X$11 VDD VSS FB 10 INVX1
X$12 VDD VSS OUT FB INVX1
.ENDS RINGO

.SUBCKT ND2X1 VDD VSS OUT B A 
M$1 OUT A VDD VDD LVPMOS L=0.25U W=1.5U 
M$2 VDD B OUT VDD LVPMOS L=0.25U W=1.5U 
M$3 VSS A 1 VSS LVNMOS L=0.25U W=0.95U 
M$4 1 B OUT VSS LVNMOS L=0.25U W=0.95U 
.ENDS ND2X1

.SUBCKT INVX1 VDD VSS OUT IN 
M$1 VDD IN OUT VDD LVPMOS L=0.25U W=1.5U 
M$2 VSS IN OUT VSS LVNMOS L=0.25U W=0.95U 
.ENDS INVX1
