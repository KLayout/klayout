* Extracted by KLayout

* cell RINGO
* pin B,FB
* pin A,ENABLE
* pin VDD
* pin OUT
* pin VSS
.SUBCKT RINGO 1 2 3 14 16
* net 1 B,FB
* net 2 A,ENABLE
* net 3 VDD
* net 14 OUT
* net 16 VSS
* cell instance $1 r0 *1 22.2,0
X$1 3 14 16 3 1 16 INVX1
* cell instance $2 r0 *1 20.4,0
X$2 3 1 16 3 13 16 INVX1
* cell instance $8 r0 *1 4.2,0
X$8 3 5 16 3 4 16 INVX1
* cell instance $9 r0 *1 6,0
X$9 3 6 16 3 5 16 INVX1
* cell instance $10 r0 *1 7.8,0
X$10 3 7 16 3 6 16 INVX1
* cell instance $11 r0 *1 9.6,0
X$11 3 8 16 3 7 16 INVX1
* cell instance $12 r0 *1 11.4,0
X$12 3 9 16 3 8 16 INVX1
* cell instance $13 r0 *1 13.2,0
X$13 3 10 16 3 9 16 INVX1
* cell instance $14 r0 *1 15,0
X$14 3 11 16 3 10 16 INVX1
* cell instance $15 r0 *1 16.8,0
X$15 3 12 16 3 11 16 INVX1
* cell instance $16 r0 *1 18.6,0
X$16 3 13 16 3 12 16 INVX1
* device instance $1 r0 *1 2.65,5.8 PMOS
M$1 3 2 4 3 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 r0 *1 3.35,5.8 PMOS
M$2 4 1 3 3 PMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 r0 *1 2.65,2.135 NMOS
M$3 15 2 16 16 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U PD=1.4U
* device instance $4 r0 *1 3.35,2.135 NMOS
M$4 4 1 15 16 NMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
.ENDS RINGO

* cell INVX1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin IN
* pin SUBSTRATE
.SUBCKT INVX1 1 2 3 4 5 6
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 IN
* net 6 SUBSTRATE
* device instance $1 r0 *1 0.85,2.135 NMOS
M$1 2 5 3 6 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $2 r0 *1 0.85,5.8 PMOS
M$2 2 5 1 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
.ENDS INVX1
