
* Simple CMOS inverer circuit 

.SUBCKT INVERTER VSS IN OUT NWELL SUBSTRATE VDD 
Mp VDD IN OUT NWELL PMOS W=1.5U L=0.25U
Mn OUT IN VSS SUBSTRATE NMOS W=0.9U L=0.25U
.ENDS

