* Extracted by KLayout

.SUBCKT TOP A Q VDD SUBSTRATE|VSS
X$1 Q SUBSTRATE|VSS VDD \$1 INV
X$2 \$1 SUBSTRATE|VSS VDD A INV
.ENDS TOP

.SUBCKT INV \$1 SUBSTRATE \$4 \$6
M$1 \$4 \$6 \$1 \$4 PMOS L=0.25U W=0.95U AS=1.02125P AD=0.73625P PS=4.05U
+ PD=3.45U
M$2 SUBSTRATE \$6 \$1 SUBSTRATE NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P
+ PS=3.45U PD=3.45U
.ENDS INV
