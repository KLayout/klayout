.subckt RINGO 11 12 13 14 15
  x$1 12 1 15 12 11 14 15 ND2X1
  x$2 12 2 15 12 1 15 INVX1
  x$3 12 3 15 12 2 15 INVX1
  x$4 12 4 15 12 3 15 INVX1
  x$5 12 5 15 12 4 15 INVX1
  x$6 12 6 15 12 5 15 INVX1
  x$7 12 7 15 12 6 15 INVX1
  x$8 12 8 15 12 7 15 INVX1
  x$9 12 9 15 12 8 15 INVX1
  x$10 12 10 15 12 9 15 INVX1
  x$11 12 11 15 12 10 15 INVX1
  x$12 12 13 15 12 11 15 INVX1
.ends RINGO

