magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 432 432 540
rect 0 216 432 324
<< properties >>
string FIXED_BBOX 0 -216 540 756
<< end >>
