magic
tech scmos
timestamp 1534318840
<< silk >>
rect 0 14 12 18
rect 4 0 8 14
<< end >>
