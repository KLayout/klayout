* Extracted by KLayout

.SUBCKT TOP
X$2 \$1 \$I2 \$I1 \$I1 \$1.Q \$2 INV2
X$3 \$1.A \$I3 \$2 \$I3 \$I2 \$1 INVCHAIN
.ENDS TOP

.SUBCKT INVCHAIN IN IN2 VSS|VSS2|VSS2B OUT OUT2 VDD
X$1 VDD IN2 \$1 \$1 OUT2 VSS|VSS2|VSS2B INV2
X$2 VDD IN \$2 \$2 OUT VSS|VSS2|VSS2B INV2
.ENDS INVCHAIN

.SUBCKT INV2 VDD A1 A2 Q1 Q2 VSS
X$1 VSS VDD A2 Q2 INV
X$2 VSS VDD A1 Q1 INV
.ENDS INV2

.SUBCKT INV \$1 \$2 \$3 \$4
M$1 \$2 \$3 \$4 \$4 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
M$2 \$1 \$3 \$4 \$4 NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
.ENDS INV
