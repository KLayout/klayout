* VDIV netlist before simplification

* cell TOP
.SUBCKT TOP 1 2 4 7
* net 1 OUT
* net 2 GND
* net 4 IN
* net 7 VDD
* device instance $1 1.025,0.335 RES, model M1
R$1 6 1 7650 M1
* device instance $2 2.85,0.335 RES, model M2
R$2 3 1 7650 M2
* device instance $3 4.665,0.335 RES, model M3
R$3 3 2 2670 M3
* device instance $4 1.765,7.485 HVPMOS
M$4 7 4 6 7 MHVPMOS L=0.25U W=1.5U AS=0.63P AD=0.63P PS=3.84U PD=3.84U
.ENDS TOP
