magic
tech scmos
timestamp 1534325915
<< silk >>
rect 0 0 12 4
<< end >>
