
* cell INVCHAIN
.SUBCKT INVCHAIN
X$2 1 2 3 4 4 5 INV2
.ENDS INVCHAIN

* cell INV2
.SUBCKT INV2 VDD VSS A1 Q1 A2 Q2 
X$1 VDD VSS A1 Q1 INV
X$2 VDD VSS A2 Q2 INV
.ENDS INV2

* cell INV
.SUBCKT INV VDD VSS A Q 
M$1 VDD A Q VDD PMOS L=0.25U W=0.95U
M$3 VSS A Q VSS NMOS L=0.25U W=0.95U
.ENDS INV

