magic
tech scmos
timestamp 1534323117
<< silk >>
rect 0 16 3 18
rect 0 14 4 16
rect 0 12 5 14
rect 8 12 12 18
rect 0 8 12 12
rect 0 0 4 8
rect 7 4 12 8
rect 8 2 12 4
rect 9 0 12 2
<< end >>
