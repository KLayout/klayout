VERSION 5.4 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
NOWIREEXTENSIONATPIN OFF ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

NONDEFAULTRULE DOUBLESPACE
    LAYER M1
        WIDTH 0.16 ;
        SPACING 0.36 ;
    END M1

# klayout 0.28.5 lef reader get's confused by the SPACING in NONDEFAULTRULE
    SPACING 
        SAMENET M1 M1 0.36 ;
    END SPACING 

END DOUBLESPACE
END LIBRARY

