magic
tech scmos
timestamp 1542205474
<< polysilicon >>
rect 130 176 170 199
rect 130 102 170 125
<< metal1 >>
rect 100 225 200 245
rect 130 219 170 225
rect 130 75 170 82
rect 100 55 200 75
<< rnfet >>
rect 130 153 170 176
<< rpfet >>
rect 130 125 170 148
<< rpoly >>
rect 130 148 170 153
<< polycontact >>
rect 130 199 170 219
rect 130 82 170 102
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_k  L500_CHAR_k_0
timestamp 1534322894
transform 1 0 145 0 1 260
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 225 0 1 140
box 0 0 12 18
use Library/magic/L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 244 0 1 151
box 0 0 16 18
use Library/magic/L500_CHAR_4  L500_CHAR_4_0
timestamp 1534324708
transform 1 0 264 0 1 151
box 0 0 12 18
use Library/magic/L500_CHAR_0  L500_CHAR_0_0
timestamp 1534325425
transform 1 0 280 0 1 151
box 0 0 12 18
use Library/magic/L500_CHAR_slash  L500_CHAR_slash_0
timestamp 1534532558
transform 1 0 296 0 1 151
box 0 0 8 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 244 0 1 129
box 0 0 12 18
use Library/magic/L500_CHAR_5  L500_CHAR_5_1
timestamp 1534324893
transform 1 0 260 0 1 129
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 145 0 1 20
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
