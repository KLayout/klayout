magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 324 108 756
rect 0 -216 108 216
<< properties >>
string FIXED_BBOX 0 -216 216 756
<< end >>
