magic
tech scmos
timestamp 1541937549
<< error_s >>
rect 10 62 14 68
rect 20 62 24 68
<< nwell >>
rect -16 80 52 92
rect -16 39 -4 80
rect 40 39 52 80
rect -16 27 52 39
<< polysilicon >>
rect 31 63 37 64
rect 31 61 32 63
rect 17 58 20 61
rect 28 59 32 61
rect 36 59 37 63
rect 28 58 37 59
<< ndiffusion >>
rect 20 67 28 68
rect 20 63 21 67
rect 27 63 28 67
rect 20 61 28 63
rect 20 56 28 58
rect 20 52 21 56
rect 27 52 28 56
rect 20 51 28 52
<< pdiffusion >>
rect 8 67 14 68
rect 8 63 9 67
rect 13 63 14 67
rect 8 62 14 63
<< metal1 >>
rect -21 108 28 116
rect -40 67 14 68
rect -40 63 9 67
rect 13 63 14 67
rect -40 62 14 63
rect 20 67 28 108
rect 20 63 21 67
rect 27 63 28 67
rect 80 64 86 103
rect 20 62 28 63
rect 31 63 86 64
rect -40 3 -34 62
rect 31 59 32 63
rect 36 59 86 63
rect 31 58 86 59
rect 20 56 28 57
rect 20 52 21 56
rect 27 52 28 56
rect 20 -3 28 52
rect 20 -11 80 -3
<< ntransistor >>
rect 20 58 28 61
<< nwpbase >>
rect -4 39 40 80
<< polycontact >>
rect 32 59 36 63
<< ndcontact >>
rect 21 63 27 67
rect 21 52 27 56
<< pdcontact >>
rect 9 63 13 67
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 -120 0 1 103
box 0 0 100 100
use L500_CHAR_s  L500_CHAR_s_0
timestamp 1534323853
transform 1 0 -19 0 1 148
box 0 0 12 18
use L500_CHAR_g  L500_CHAR_g_0
timestamp 1534322005
transform 1 0 64 0 1 147
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 80 0 1 103
box 0 0 100 100
use L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 98 0 1 79
box 0 0 8 18
use L500_CHAR_s  L500_CHAR_s_1
timestamp 1534323853
transform 1 0 108 0 1 79
box 0 0 12 18
use L500_CHAR_o  L500_CHAR_o_0
timestamp 1534323159
transform 1 0 122 0 1 79
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 137 0 1 79
box 0 0 12 18
use L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 97 0 1 58
box 0 0 16 18
use L500_CHAR_4  L500_CHAR_4_0
timestamp 1534324830
transform 1 0 116 0 1 58
box 0 0 12 18
use L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 97 0 1 36
box 0 0 12 18
use L500_CHAR_1  L500_CHAR_1_1
timestamp 1534326485
transform 1 0 112 0 1 36
box 0 0 12 18
use L500_CHAR_dot  L500_CHAR_dot_1
timestamp 1534325697
transform 1 0 126 0 1 36
box 0 0 4 4
use L500_CHAR_5  L500_CHAR_5_1
timestamp 1534324893
transform 1 0 132 0 1 36
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 -120 0 1 -97
box 0 0 100 100
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 -16 0 1 -61
box 0 0 12 18
use L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 64 0 1 -65
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 80 0 1 -97
box 0 0 100 100
<< end >>
