* Extracted by KLayout

* cell top
* pin FB
* pin VDD
* pin OUT
* pin ENABLE
* pin VSS
.SUBCKT top 11 12 13 14 15
* net 11 FB
* net 12 VDD
* net 13 OUT
* net 14 ENABLE
* net 15 VSS
* cell instance $1 r0 *1 1.8,0
X$1 12 1 15 12 11 14 15 nd2X1
* cell instance $2 r0 *1 4.2,0
X$2 12 2 15 12 1 15 INV
* cell instance $3 r0 *1 6,0
X$3 12 3 15 12 2 15 INV
* cell instance $4 r0 *1 7.8,0
X$4 12 4 15 12 3 15 INV
* cell instance $5 r0 *1 9.6,0
X$5 12 5 15 12 4 15 INV
* cell instance $6 r0 *1 11.4,0
X$6 12 6 15 12 5 15 INV
* cell instance $7 r0 *1 13.2,0
X$7 12 7 15 12 6 15 INV
* cell instance $8 r0 *1 15,0
X$8 12 8 15 12 7 15 INV
* cell instance $9 r0 *1 16.8,0
X$9 12 9 15 12 8 15 INV
* cell instance $10 r0 *1 18.6,0
X$10 12 10 15 12 9 15 INV
* cell instance $11 r0 *1 20.4,0
X$11 12 11 15 12 10 15 INV
* cell instance $12 r0 *1 22.2,0
X$12 12 13 15 12 11 15 INV
.ENDS top

* cell INV
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin IN
* pin SUBSTRATE
.SUBCKT INV 1 2 3 4 5 6
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 IN
* net 6 SUBSTRATE
* device instance $1 r0 *1 0.85,5.8 PMOS
M$1 2 5 1 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $2 r0 *1 0.85,2.135 NMOS
M$2 2 5 3 6 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
.ENDS INV

* cell nd2X1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin B
* pin A
* pin SUBSTRATE
.SUBCKT nd2X1 1 2 3 4 5 6 7
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 B
* net 6 A
* net 7 SUBSTRATE
* device instance $1 r0 *1 0.85,5.8 PMOS
M$1 1 6 2 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 r0 *1 1.55,5.8 PMOS
M$2 2 5 1 4 PMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 r0 *1 0.85,2.135 NMOS
M$3 8 6 3 7 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U PD=1.4U
* device instance $4 r0 *1 1.55,2.135 NMOS
M$4 2 5 8 7 NMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
.ENDS nd2X1
