VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.05 ;

LAYER M1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  WIDTH		0.2 ;
END M1

LAYER V2
  TYPE	CUT ;
END V2

LAYER M2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  WIDTH		0.2 ;
END M2

VIA M2_M1 DEFAULT
  LAYER M1 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER V2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER M2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END M2_M1

END LIBRARY
