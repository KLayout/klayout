magic
tech scmos
timestamp 1533916061
<< pwell >>
rect 6 404 334 436
rect 404 274 436 594
<< nwell >>
rect 164 6 196 326
rect 274 164 594 196
<< polysilicon >>
rect 419 584 421 586
rect 14 419 16 421
rect 324 419 335 421
rect 179 316 181 327
rect 419 273 421 284
rect 273 179 284 181
rect 584 179 586 181
rect 179 14 181 16
<< ndiffusion >>
rect 20 422 320 426
rect 16 421 324 422
rect 16 418 324 419
rect 20 414 320 418
rect 418 580 419 584
rect 414 288 419 580
rect 418 284 419 288
rect 421 580 422 584
rect 421 288 426 580
rect 421 284 422 288
<< pdiffusion >>
rect 178 312 179 316
rect 174 20 179 312
rect 178 16 179 20
rect 181 312 182 316
rect 181 20 186 312
rect 181 16 182 20
rect 288 182 580 186
rect 284 181 584 182
rect 284 178 584 179
rect 288 174 580 178
<< metal1 >>
rect 352 588 418 592
rect 414 584 418 588
rect 8 426 12 500
rect 328 426 332 430
rect 8 422 16 426
rect 324 422 332 426
rect 336 422 340 488
rect 328 418 332 422
rect 339 418 340 422
rect 8 414 16 418
rect 324 414 332 418
rect 8 352 12 414
rect 328 410 332 414
rect 328 352 332 406
rect 112 331 182 332
rect 112 328 178 331
rect 170 320 190 324
rect 174 316 178 320
rect 182 316 186 320
rect 174 12 178 16
rect 112 8 178 12
rect 194 320 248 324
rect 352 276 406 280
rect 422 588 488 592
rect 422 584 426 588
rect 414 280 418 284
rect 422 280 426 284
rect 410 276 430 280
rect 422 269 488 272
rect 418 268 488 269
rect 276 194 280 248
rect 276 186 280 190
rect 588 186 592 248
rect 276 182 284 186
rect 584 182 592 186
rect 269 112 273 178
rect 276 178 280 182
rect 276 174 284 178
rect 584 174 592 178
rect 276 170 280 174
rect 588 112 592 174
rect 182 12 186 16
rect 182 8 248 12
<< ntransistor >>
rect 16 419 324 421
rect 419 284 421 584
<< ptransistor >>
rect 179 16 181 316
rect 284 179 584 181
<< polycontact >>
rect 335 418 339 422
rect 178 327 182 331
rect 418 269 422 273
rect 269 178 273 182
<< ndcontact >>
rect 16 422 20 426
rect 320 422 324 426
rect 16 414 20 418
rect 320 414 324 418
rect 414 580 418 584
rect 414 284 418 288
rect 422 580 426 584
rect 422 284 426 288
<< pdcontact >>
rect 174 312 178 316
rect 174 16 178 20
rect 182 312 186 316
rect 182 16 186 20
rect 284 182 288 186
rect 580 182 584 186
rect 284 174 288 178
rect 580 174 584 178
<< psubstratepcontact >>
rect 16 430 332 434
rect 16 406 332 410
rect 406 276 410 584
rect 430 276 434 584
<< nsubstratencontact >>
rect 166 16 170 324
rect 190 16 194 324
rect 276 190 584 194
rect 276 166 584 170
<< nplusdoping >>
rect 170 320 179 324
rect 181 320 190 324
rect 584 190 592 194
rect 276 181 280 190
rect 276 170 280 179
rect 588 170 592 190
rect 584 166 592 170
rect 166 12 170 16
rect 190 12 194 16
rect 166 8 194 12
<< pplusdoping >>
rect 406 588 434 592
rect 406 584 410 588
rect 430 584 434 588
rect 8 430 16 434
rect 8 410 12 430
rect 328 421 332 430
rect 328 410 332 419
rect 8 406 16 410
rect 410 276 419 280
rect 421 276 430 280
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_6 Library/magic
timestamp 1531942424
transform 1 0 0 0 1 480
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_7
timestamp 1531942424
transform 1 0 240 0 1 480
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_8
timestamp 1531942424
transform 1 0 480 0 1 480
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_1
timestamp 1531942424
transform 1 0 0 0 1 240
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_3
timestamp 1531942424
transform 1 0 240 0 1 240
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_5
timestamp 1531942424
transform 1 0 480 0 1 240
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_0
timestamp 1531942424
transform 1 0 0 0 1 0
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_2
timestamp 1531942424
transform 1 0 240 0 1 0
box 0 0 120 120
use Library/magic/L500_TPM1_blank  L500_TPM1_blank_4
timestamp 1531942424
transform 1 0 480 0 1 0
box 0 0 120 120
<< labels >>
rlabel space 260 260 340 340 1 gnd!
rlabel space 20 500 100 580 1 DRAIN_NMOS0
rlabel space 500 500 580 580 1 DRAIN_NMOS1
rlabel space 500 20 580 100 1 DRAIN_PMOS0
rlabel space 20 20 100 100 1 DRAIN_PMOS0
rlabel space 260 500 340 580 1 GATE_NMOS0
rlabel space 500 260 580 340 1 GATE_NMOS1
rlabel space 260 20 340 100 1 GATE_PMOS0
rlabel space 20 260 100 340 1 GATE_PMOS1
<< end >>
