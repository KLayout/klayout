
.SUBCKT RINGO VSS VDD FB ENABLE OUT
X$1 VDD 1 VSS VDD FB ENABLE VSS ND2X1
X$2 VDD 2 VSS VDD 1 VSS INVX1
X$3 VDD 3 VSS VDD 2 VSS INVX1
X$4 VDD 4 VSS VDD 3 VSS INVX1
X$5 VDD 5 VSS VDD 4 VSS INVX1
X$6 VDD 6 VSS VDD 5 VSS INVX1
X$7 VDD 7 VSS VDD 6 VSS INVX1
X$8 VDD 8 VSS VDD 7 VSS INVX1
X$9 VDD 9 VSS VDD 8 VSS INVX1
X$10 VDD 10 VSS VDD 9 VSS INVX1
X$11 VDD FB VSS VDD 10 VSS INVX1
X$12 VDD OUT VSS VDD FB VSS INVX1
.ENDS RINGO

.SUBCKT ND2X1 VDD OUT VSS NWELL B A BULK
M$1 OUT A VDD NWELL PMOS L=0.251U W=1.6U 
M$2 VDD B OUT NWELL PMOS L=0.25U W=1.5U 
M$3 VSS A 1 BULK NMOS L=0.26U W=1.00U 
M$4 1 B OUT BULK NMOS L=0.25U W=0.95U 
.ENDS ND2X1

.SUBCKT INVX1 VDD OUT VSS NWELL IN BULK
M$1 VDD IN OUT NWELL PMOS L=0.25U W=1.5U 
M$2 VSS IN OUT BULK NMOS L=0.25U W=0.95U 
.ENDS INVX1
