LAYER OD
    TYPE IMPLANT ;
END OD
LAYER VTS_N
    TYPE IMPLANT ;
END VTS_N
LAYER VTS_P
    TYPE IMPLANT ;
END VTS_P
LAYER M0OD
    TYPE IMPLANT ;
END M0OD
LAYER M0PO 
    TYPE MASTERSLICE ;
END M0PO
LAYER VIA0
    TYPE CUT ;
END VIA0
LAYER M1
    TYPE MASTERSLICE ;
END M1
LAYER VIA1
    TYPE CUT ;
END VIA1
LAYER M2
    TYPE MASTERSLICE ;
END M2

VIA square 
    LAYER M0PO ;
        RECT -0.006 -0.006 0.006 0.006 ;
    LAYER VIA0 ;
        RECT -0.006 -0.006 0.006 0.006 ;
    LAYER M1 ;
        RECT -0.006 -0.006 0.006 0.006 ;
END square
