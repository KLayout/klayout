* Extracted by KLayout

.SUBCKT INVCHAIN IN OUT VSS VDD
X$1 IN \$2 \$3 \$2 \$3 \$4 VDD VSS INV3
X$2 \$5 \$6 \$4 \$5 VDD VSS INV2
X$3 VSS VDD \$6 OUT INV
.ENDS INVCHAIN

.SUBCKT INV2 \$I8 \$I7 \$I6 \$I5 \$I4 \$I2
X$1 \$I2 \$I4 \$I6 \$I8 INV
X$2 \$I2 \$I4 \$I5 \$I7 INV
.ENDS INV2

.SUBCKT INV3 3 5 7 4 6 8 \$I4 \$I2
X$1 \$I2 \$I4 3 4 INV
X$2 \$I2 \$I4 5 6 INV
X$3 \$I2 \$I4 7 8 INV
.ENDS INV3

.SUBCKT INV \$1 \$2 \$3 \$4
M$1 \$2 \$3 \$4 \$4 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.5225P PS=3.45U PD=3U
M$2 \$1 \$3 \$4 \$4 NMOS L=0.25U W=0.95U AS=0.73625P AD=0.5225P PS=3.45U PD=3U
.ENDS INV
