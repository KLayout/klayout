magic
tech scmos
timestamp 1534321786
<< silk >>
rect 1 16 12 18
rect 0 15 12 16
rect 0 12 4 15
rect 0 8 12 12
rect 0 5 4 8
rect 0 4 5 5
rect 0 2 12 4
rect 2 0 12 2
<< end >>
