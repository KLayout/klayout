* Extracted by KLayout

.SUBCKT INVCHAIN ANY R ANY$1 PWR GND
X$1 ANY R R ANY$1 PWR GND INV2
.ENDS INVCHAIN

.SUBCKT INV2 A1 A2 Q1 Q2 R VSS
X$1 VSS R A1 Q1 INV
X$2 VSS R A2 Q2 INV
.ENDS INV2

.SUBCKT INV \$1 \$2 \$3 \$4
M$1 \$2 \$3 \$4 \$4 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
M$2 \$1 \$3 \$4 \$4 NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
.ENDS INV
