magic
tech scmos
timestamp 1538327581
<< polysilicon >>
rect 111 75 903 83
<< metal1 >>
rect 100 75 103 83
rect 911 75 914 83
<< polycontact >>
rect 103 75 111 83
rect 903 75 911 83
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 914 0 1 0
box 0 0 100 100
<< end >>
