LAYER M0PO 
    TYPE MASTERSLICE ;
    WIDTH 0.02 ;
END M0PO
LAYER VIA0
    TYPE CUT ;
END VIA0
LAYER M1
    TYPE MASTERSLICE ;
    WIDTH 0.025 ;
END M1
LAYER VIA1
    TYPE CUT ;
END VIA1
LAYER M2
    TYPE MASTERSLICE ;
    WIDTH 0.03 ;
END M2

VIA square 
    LAYER M0PO ;
        RECT -0.006 -0.006 0.006 0.006 ;
    LAYER VIA0 ;
        RECT -0.006 -0.006 0.006 0.006 ;
    LAYER M1 ;
        RECT -0.006 -0.006 0.006 0.006 ;
END square
