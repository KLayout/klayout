magic
tech scmos
timestamp 1534532558
<< silk >>
rect 4 15 8 18
rect 3 14 8 15
rect 3 11 7 14
rect 2 7 6 11
rect 1 4 5 7
rect 0 3 5 4
rect 0 0 4 3
<< end >>
