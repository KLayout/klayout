VERSION 5.7 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO POLYGON_PIN
  FOREIGN POLYGON_PIN ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 200.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        POLYGON 0.000 10.000 30.000 10.000 30.000 0.000 35.000 0.000 35.000 15.000 0.000 15.0000 ;
    END
  END VDD
END POLYGON_PIN

END LIBRARY

