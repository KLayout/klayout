magic
tech scmos
timestamp 1538315839
<< metal1 >>
rect 108 280 200 285
rect 108 192 192 280
rect 280 192 285 200
rect 15 108 285 192
rect 15 100 20 108
rect 108 20 192 108
rect 100 15 192 20
<< metal2 >>
rect 100 280 192 285
rect 15 192 20 200
rect 108 192 192 280
rect 15 108 285 192
rect 108 20 192 108
rect 280 100 285 108
rect 108 15 200 20
use Library/magic/L500_CHAR_m  L500_CHAR_m_0 Library/magic
timestamp 1534323034
transform 1 0 4 0 1 304
box 0 0 16 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0 Library/magic
timestamp 1534321786
transform 1 0 24 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_t  L500_CHAR_t_0 Library/magic
timestamp 1534318840
transform 1 0 40 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0 Library/magic
timestamp 1534325357
transform 1 0 56 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_0 Library/magic
timestamp 1534225390
transform 1 0 72 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_0 Library/magic
timestamp 1534324708
transform 1 0 88 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_slash  L500_CHAR_slash_0 Library/magic
timestamp 1534532558
transform 1 0 104 0 1 304
box 0 0 8 18
use Library/magic/L500_CHAR_m  L500_CHAR_m_1
timestamp 1534323034
transform 1 0 116 0 1 304
box 0 0 16 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_1
timestamp 1534321786
transform 1 0 136 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_t  L500_CHAR_t_1
timestamp 1534318840
transform 1 0 152 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_1
timestamp 1534325357
transform 1 0 168 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_1
timestamp 1534225390
transform 1 0 184 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_0 Library/magic
timestamp 1534326485
transform 1 0 200 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_under  L500_CHAR_under_0 Library/magic
timestamp 1534325915
transform 1 0 216 0 1 304
box 0 0 12 4
use Library/magic/L500_CHAR_c  L500_CHAR_c_0 Library/magic
timestamp 1534321654
transform 1 0 232 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_2
timestamp 1534325357
transform 1 0 248 0 1 304
box 0 0 12 18
use Library/magic/L500_CHAR_p  L500_CHAR_p_0 Library/magic
timestamp 1534323210
transform 1 0 264 0 1 304
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2 Library/magic
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
