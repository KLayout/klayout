
.SUBCKT NAND2_WITH_DIODES A B OUT VSS VDD
M1 VDD B OUT VDD PMOS L=0.25U W=1.5U
M2 VDD A OUT VDD PMOS L=0.25U W=1.5U
M3 VSS B $1 VSS NMOS L=0.25U W=1.8U
M4 $1 A OUT VSS NMOS L=0.25U W=1.8U
.ENDS 
