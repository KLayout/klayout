* RINGO netlist

* cell RINGO
.SUBCKT RINGO
* net 1 FB
* net 2 OSC
* net 3 NEXT
* net 4 VSSZ,VSS
* net 5 VDDZ,VDD
* cell instance $1 r180 *1 -0.24,9.18
X$1 16 1 2 4 5 INV2
* cell instance $2 r0 *1 0,0
X$2 1 14 15 4 5 INV2
* cell instance $3 r180 *1 10.32,9.18
X$3 3 9 19 4 5 INV2
* cell instance $4 r0 *1 10.56,0
X$4 20 10 3 4 5 INV2
* cell instance $5 r180 *1 7.68,9.18
X$5 19 8 18 4 5 INV2
* cell instance $6 r180 *1 5.04,9.18
X$6 18 7 17 4 5 INV2
* cell instance $7 r180 *1 2.4,9.18
X$7 17 6 16 4 5 INV2
* cell instance $8 r0 *1 2.64,0
X$8 15 13 22 4 5 INV2
* cell instance $9 r0 *1 5.28,0
X$9 22 12 21 4 5 INV2
* cell instance $10 r0 *1 7.92,0
X$10 21 11 20 4 5 INV2
.ENDS RINGO

* cell INV2
* pin IN
* pin 
* pin OUT
* pin 
* pin 
.SUBCKT INV2 1 2 3 4 5
* net 1 IN
* net 3 OUT
* cell instance $1 r0 *1 -0.4,0
X$1 2 4 1 TRANS
* cell instance $2 r0 *1 -0.4,2.8
X$2 2 5 1 TRANS
* cell instance $3 m0 *1 0.4,2.8
X$3 5 3 2 TRANS
* cell instance $4 m0 *1 0.4,0
X$4 4 3 2 TRANS
* device instance $1 -0.4,0 PMOS
M$1 2 1 4 2 PMOS L=0.25U W=0.95U AS=0.49875P AD=0.26125P PS=2.95U PD=1.5U
* device instance $2 0.4,0 PMOS
M$2 4 2 3 4 PMOS L=0.25U W=0.95U AS=0.26125P AD=0.49875P PS=1.5U PD=2.95U
* device instance $3 -0.4,2.8 PMOS
M$3 2 1 5 2 PMOS L=0.25U W=0.95U AS=0.49875P AD=0.26125P PS=2.95U PD=1.5U
* device instance $4 0.4,2.8 PMOS
M$4 5 2 3 5 PMOS L=0.25U W=0.95U AS=0.26125P AD=0.49875P PS=1.5U PD=2.95U
* device instance $5 -0.4,0 NMOS
M$5 2 1 4 2 NMOS L=0.25U W=0.95U AS=0.49875P AD=0.26125P PS=2.95U PD=1.5U
* device instance $6 0.4,0 NMOS
M$6 4 2 3 4 NMOS L=0.25U W=0.95U AS=0.26125P AD=0.49875P PS=1.5U PD=2.95U
.ENDS INV2

* cell TRANS
* pin 
* pin 
* pin 
.SUBCKT TRANS 1 2 3
.ENDS TRANS
