magic
tech scmos
timestamp 1541212842
<< silk >>
rect 0 17 3 18
rect 0 14 4 17
rect 1 12 4 14
<< end >>
