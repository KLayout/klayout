magic
tech scmos
timestamp 1534324995
<< silk >>
rect 0 17 10 18
rect 0 16 11 17
rect 0 14 12 16
rect 7 13 12 14
rect 8 0 12 13
<< end >>
