magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 72 720 252 756
rect 36 684 288 720
rect 0 612 324 684
rect 0 144 108 612
rect 216 144 324 612
rect 0 72 324 144
rect 36 36 288 72
rect 72 0 252 36
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
