.subckt top r1 r2
r5  r1 r2 50.1
.ends
