* Extracted by KLayout

.SUBCKT INVCHAIN IN OUT VSS VDD
X$1 VDD IN \$1 \$1 OUT VSS INV2
.ENDS INVCHAIN

.SUBCKT INV2 VDD A1 A2 Q1 Q2 VSS
X$1 VSS VDD A2 Q2 INV
X$2 VSS VDD A1 Q1 INV
.ENDS INV2

.SUBCKT INV \$1 \$2 \$3 \$4
M$1 \$4 \$3 \$2 \$4 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
M$2 \$4 \$3 \$1 \$4 NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
.ENDS INV
