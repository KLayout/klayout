magic
tech scmos
timestamp 1534322894
<< silk >>
rect 0 11 4 18
rect 8 15 12 18
rect 7 13 12 15
rect 7 11 11 13
rect 0 7 10 11
rect 0 0 4 7
rect 7 5 11 7
rect 7 3 12 5
rect 8 0 12 3
<< end >>
