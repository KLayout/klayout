magic
tech scmos
timestamp 1542451143
<< nwell >>
rect 113 178 187 188
rect 113 141 123 178
rect 177 141 187 178
rect 113 129 187 141
<< metal1 >>
rect 100 200 139 210
rect 129 173 139 200
rect 161 200 200 210
rect 161 173 171 200
rect 129 165 171 173
rect 129 147 135 165
rect 165 163 171 165
rect 138 156 162 162
rect 138 100 144 156
rect 100 90 144 100
rect 147 152 153 153
rect 147 148 148 152
rect 152 148 153 152
rect 147 100 153 148
rect 156 147 162 156
rect 165 148 166 163
rect 170 148 171 163
rect 165 147 171 148
rect 147 90 200 100
<< nwpbase >>
rect 123 173 177 178
rect 123 146 128 173
rect 136 154 164 164
rect 136 146 146 154
rect 154 146 164 154
rect 172 146 177 173
rect 123 145 147 146
rect 153 145 177 146
rect 123 141 177 145
<< nwpnbase >>
rect 128 164 172 173
rect 128 146 136 164
rect 146 146 154 154
rect 164 146 172 164
rect 147 145 153 146
<< pbasepdiffcontact >>
rect 139 157 161 161
rect 139 148 143 157
rect 157 148 161 157
<< nbasendiffcontact >>
rect 130 167 170 171
rect 130 148 134 163
<< ndcontact >>
rect 148 148 152 152
rect 166 148 170 163
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_c  L500_CHAR_c_0
timestamp 1534321654
transform 1 0 136 0 1 232
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 199 0 1 169
box 0 0 12 18
use Library/magic/L500_CHAR_p  L500_CHAR_p_0
timestamp 1534323210
transform 1 0 215 0 1 169
box 0 0 12 18
use Library/magic/L500_CHAR_n  L500_CHAR_n_1
timestamp 1534323117
transform 1 0 231 0 1 169
box 0 0 12 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_0
timestamp 1534324708
transform 1 0 247 0 1 169
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 199 0 1 147
box 0 0 8 18
use Library/magic/L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 32 0 1 113
box 0 0 12 18
use Library/magic/L500_CHAR_e  L500_CHAR_e_0
timestamp 1534321786
transform 1 0 209 0 1 109
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
