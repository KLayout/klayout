* Extracted by KLayout

* cell SP6TArray_2X4
.SUBCKT SP6TArray_2X4
* net 1 vdd
* net 2 bl[0]
* net 3 bl_n[0]
* net 4 bl[1]
* net 5 bl_n[1]
* net 6 bl[2]
* net 7 bl_n[2]
* net 8 bl[3]
* net 9 bl_n[3]
* net 26 wl[0]
* net 31 wl[1]
* net 52 vss
* device instance $1 r0 *1 0.215,1.935 sky130_fd_pr__nfet_01v8__model
M$1 52 11 12 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.1113P
+ AD=0.18165P PS=1.37U PD=1.285U
* device instance $2 r0 *1 0.605,2.56 sky130_fd_pr__nfet_01v8__model
M$2 12 26 2 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $3 r0 *1 0.605,2.99 sky130_fd_pr__nfet_01v8__model
M$3 2 31 32 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $4 r0 *1 0.215,3.615 sky130_fd_pr__nfet_01v8__model
M$4 32 34 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.1113P PS=1.285U PD=1.37U
* device instance $5 r0 *1 1.965,1.935 sky130_fd_pr__nfet_01v8__model
M$5 11 12 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $6 r0 *1 2.395,1.935 sky130_fd_pr__nfet_01v8__model
M$6 52 15 16 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $7 r0 *1 1.575,2.56 sky130_fd_pr__nfet_01v8__model
M$7 11 26 3 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $8 r0 *1 2.785,2.56 sky130_fd_pr__nfet_01v8__model
M$8 16 26 4 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $9 r0 *1 1.575,2.99 sky130_fd_pr__nfet_01v8__model
M$9 3 31 34 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $10 r0 *1 2.785,2.99 sky130_fd_pr__nfet_01v8__model
M$10 4 31 35 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $11 r0 *1 1.965,3.615 sky130_fd_pr__nfet_01v8__model
M$11 34 32 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $12 r0 *1 2.395,3.615 sky130_fd_pr__nfet_01v8__model
M$12 35 37 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $13 r0 *1 4.145,1.935 sky130_fd_pr__nfet_01v8__model
M$13 15 16 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $14 r0 *1 4.575,1.935 sky130_fd_pr__nfet_01v8__model
M$14 52 19 20 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $15 r0 *1 3.755,2.56 sky130_fd_pr__nfet_01v8__model
M$15 15 26 5 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $16 r0 *1 4.965,2.56 sky130_fd_pr__nfet_01v8__model
M$16 20 26 6 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $17 r0 *1 3.755,2.99 sky130_fd_pr__nfet_01v8__model
M$17 5 31 37 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $18 r0 *1 4.965,2.99 sky130_fd_pr__nfet_01v8__model
M$18 6 31 38 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $19 r0 *1 4.145,3.615 sky130_fd_pr__nfet_01v8__model
M$19 37 35 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $20 r0 *1 4.575,3.615 sky130_fd_pr__nfet_01v8__model
M$20 38 40 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $21 r0 *1 6.325,1.935 sky130_fd_pr__nfet_01v8__model
M$21 19 20 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $22 r0 *1 6.755,1.935 sky130_fd_pr__nfet_01v8__model
M$22 52 23 24 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $23 r0 *1 5.935,2.56 sky130_fd_pr__nfet_01v8__model
M$23 19 26 7 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $24 r0 *1 7.145,2.56 sky130_fd_pr__nfet_01v8__model
M$24 24 26 8 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $25 r0 *1 5.935,2.99 sky130_fd_pr__nfet_01v8__model
M$25 7 31 40 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $26 r0 *1 7.145,2.99 sky130_fd_pr__nfet_01v8__model
M$26 8 31 41 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $27 r0 *1 6.325,3.615 sky130_fd_pr__nfet_01v8__model
M$27 40 38 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $28 r0 *1 6.755,3.615 sky130_fd_pr__nfet_01v8__model
M$28 41 50 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $29 r0 *1 8.505,1.935 sky130_fd_pr__nfet_01v8__model
M$29 23 24 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.1113P PS=1.285U PD=1.37U
* device instance $30 r0 *1 8.115,2.56 sky130_fd_pr__nfet_01v8__model
M$30 23 26 9 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.0588P PS=1.285U PD=0.7U
* device instance $31 r0 *1 8.115,2.99 sky130_fd_pr__nfet_01v8__model
M$31 9 31 50 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.18165P PS=0.7U PD=1.285U
* device instance $32 r0 *1 8.505,3.615 sky130_fd_pr__nfet_01v8__model
M$32 50 41 52 52 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.1113P PS=1.285U PD=1.37U
* device instance $33 r0 *1 0.215,0.605 sky130_fd_pr__pfet_01v8__model
M$33 1 11 12 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1113P
+ AD=0.1869P PS=1.37U PD=1.73U
* device instance $34 r0 *1 1.965,0.605 sky130_fd_pr__pfet_01v8__model
M$34 11 12 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.0588P PS=1.73U PD=0.7U
* device instance $35 r0 *1 2.395,0.605 sky130_fd_pr__pfet_01v8__model
M$35 1 15 16 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.1869P PS=0.7U PD=1.73U
* device instance $36 r0 *1 4.145,0.605 sky130_fd_pr__pfet_01v8__model
M$36 15 16 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.0588P PS=1.73U PD=0.7U
* device instance $37 r0 *1 4.575,0.605 sky130_fd_pr__pfet_01v8__model
M$37 1 19 20 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.1869P PS=0.7U PD=1.73U
* device instance $38 r0 *1 6.325,0.605 sky130_fd_pr__pfet_01v8__model
M$38 19 20 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.0588P PS=1.73U PD=0.7U
* device instance $39 r0 *1 6.755,0.605 sky130_fd_pr__pfet_01v8__model
M$39 1 23 24 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.1869P PS=0.7U PD=1.73U
* device instance $40 r0 *1 8.505,0.605 sky130_fd_pr__pfet_01v8__model
M$40 23 24 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.1113P PS=1.73U PD=1.37U
* device instance $41 r0 *1 0.215,4.945 sky130_fd_pr__pfet_01v8__model
M$41 1 34 32 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1113P
+ AD=0.1869P PS=1.37U PD=1.73U
* device instance $42 r0 *1 1.965,4.945 sky130_fd_pr__pfet_01v8__model
M$42 34 32 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.0588P PS=1.73U PD=0.7U
* device instance $43 r0 *1 2.395,4.945 sky130_fd_pr__pfet_01v8__model
M$43 1 37 35 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.1869P PS=0.7U PD=1.73U
* device instance $44 r0 *1 4.145,4.945 sky130_fd_pr__pfet_01v8__model
M$44 37 35 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.0588P PS=1.73U PD=0.7U
* device instance $45 r0 *1 4.575,4.945 sky130_fd_pr__pfet_01v8__model
M$45 1 40 38 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.1869P PS=0.7U PD=1.73U
* device instance $46 r0 *1 6.325,4.945 sky130_fd_pr__pfet_01v8__model
M$46 40 38 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.0588P PS=1.73U PD=0.7U
* device instance $47 r0 *1 6.755,4.945 sky130_fd_pr__pfet_01v8__model
M$47 1 50 41 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.0588P
+ AD=0.1869P PS=0.7U PD=1.73U
* device instance $48 r0 *1 8.505,4.945 sky130_fd_pr__pfet_01v8__model
M$48 50 41 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.1113P PS=1.73U PD=1.37U
.ENDS SP6TArray_2X4
