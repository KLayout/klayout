magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 72 720 324 756
rect 36 684 324 720
rect 0 612 324 684
rect 0 468 108 612
rect 0 432 252 468
rect 0 396 288 432
rect 36 360 324 396
rect 72 324 324 360
rect 216 144 324 324
rect 0 72 324 144
rect 0 36 288 72
rect 0 0 252 36
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
