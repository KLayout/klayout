* Extracted by KLayout

* cell Rre
* pin gnd!
* pin vdd!
.SUBCKT Rre 1 2
* net 1 gnd!
* net 2 vdd!
* device instance $1 r0 *1 8.43,1.51 RR1
R$1 1 2 10 RR1 L=6U W=0.6U
.ENDS Rre
