* Extracted by KLayout

* cell TOP
.SUBCKT TOP
* net 1 4
* net 2 3
* net 3 2
* net 4 1
* net 5 8
* net 6 7
* net 7 5
* net 8 6
* cell instance $1 r0 *1 0,0
X$1 1 2 7 3 4 5 8 6 CHIP
.ENDS TOP

* cell CHIP
* pin pad3
* pin pad4
* pin pad5
* pin pad2
* pin pad1
* pin pad8
* pin pad6
* pin pad7
.SUBCKT CHIP 1 2 3 4 5 6 7 8
.ENDS CHIP
