magic
tech scmos
timestamp 1534324403
<< silk >>
rect 0 12 4 18
rect 8 12 12 18
rect 0 10 12 12
rect 1 9 11 10
rect 2 8 10 9
rect 3 6 9 8
rect 4 0 8 6
<< end >>
