magic
tech scmos
timestamp 1541938952
<< error_s >>
rect 11 65 15 66
rect 21 65 25 71
<< nwell >>
rect -15 83 53 95
rect -15 37 -3 83
rect 41 37 53 83
rect -15 25 53 37
<< polysilicon >>
rect 18 56 21 64
rect 29 63 38 64
rect 29 57 33 63
rect 37 57 38 63
rect 29 56 38 57
<< ndiffusion >>
rect 21 70 29 71
rect 21 66 22 70
rect 28 66 29 70
rect 21 64 29 66
rect 21 54 29 56
rect 21 50 22 54
rect 28 50 29 54
rect 21 49 29 50
<< pdiffusion >>
rect 9 70 15 71
rect 9 66 10 70
rect 14 66 15 70
rect 9 65 15 66
<< metal1 >>
rect -21 108 29 116
rect -54 70 15 71
rect -54 66 10 70
rect 14 66 15 70
rect -54 65 15 66
rect 21 70 29 108
rect 21 66 22 70
rect 28 66 29 70
rect 21 65 29 66
rect -54 2 -48 65
rect 86 64 94 103
rect 32 63 94 64
rect 32 57 33 63
rect 37 57 94 63
rect 32 56 94 57
rect 21 54 29 55
rect 21 50 22 54
rect 28 50 29 54
rect 21 -8 29 50
rect 21 -16 81 -8
<< ntransistor >>
rect 21 56 29 64
<< nwpbase >>
rect -3 37 41 83
<< polycontact >>
rect 33 57 37 63
<< ndcontact >>
rect 22 66 28 70
rect 22 50 28 54
<< pdcontact >>
rect 10 66 14 70
use L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 -120 0 1 103
box 0 0 100 100
use L500_CHAR_s  L500_CHAR_s_0
timestamp 1534323853
transform 1 0 -19 0 1 148
box 0 0 12 18
use L500_CHAR_g  L500_CHAR_g_0
timestamp 1534322005
transform 1 0 64 0 1 147
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 80 0 1 103
box 0 0 100 100
use L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 98 0 1 79
box 0 0 8 18
use L500_CHAR_s  L500_CHAR_s_1
timestamp 1534323853
transform 1 0 108 0 1 79
box 0 0 12 18
use L500_CHAR_o  L500_CHAR_o_0
timestamp 1534323159
transform 1 0 122 0 1 79
box 0 0 12 18
use L500_CHAR_n  L500_CHAR_n_0
timestamp 1534323117
transform 1 0 137 0 1 79
box 0 0 12 18
use L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 97 0 1 58
box 0 0 16 18
use L500_CHAR_4  L500_CHAR_4_0
timestamp 1534324830
transform 1 0 116 0 1 58
box 0 0 12 18
use L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 97 0 1 36
box 0 0 12 18
use L500_CHAR_4  L500_CHAR_4_1
timestamp 1534324830
transform 1 0 111 0 1 36
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 -120 0 1 -97
box 0 0 100 100
use L500_CHAR_b  L500_CHAR_b_0
timestamp 1534321628
transform 1 0 -16 0 1 -61
box 0 0 12 18
use L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 64 0 1 -65
box 0 0 12 18
use L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 80 0 1 -97
box 0 0 100 100
<< end >>
