* Extracted by KLayout

.SUBCKT TOP A Q VDD SUBSTRATE|VSS
X$1 SUBSTRATE|VSS VDD VDD \$1 Q SUBSTRATE|VSS INV
X$2 SUBSTRATE|VSS VDD VDD A \$1 SUBSTRATE|VSS INV
.ENDS TOP

.SUBCKT INV \$1 \$2 \$3 \$4 \$5 SUBSTRATE
M$1 \$2 \$4 \$5 \$3 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
M$2 \$1 \$4 \$5 SUBSTRATE NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
.ENDS INV
