* Extracted by KLayout

* cell RINGO
* pin FB
* pin VDD
* pin OUT
* pin ENABLE
* pin VSS
.SUBCKT RINGO 11 12 13 14 15
* net 11 FB
* net 12 VDD
* net 13 OUT
* net 14 ENABLE
* net 15 VSS
* cell instance $1 r0 *1 1.8,0
X$1 12 1 15 12 11 14 15 ND2X1
* cell instance $2 r0 *1 4.7,0
X$2 12 2 15 12 1 15 INVX1
* cell instance $3 r0 *1 6.5,0
X$3 12 3 15 12 2 15 INVX1
* cell instance $4 r0 *1 8.3,0
X$4 12 4 15 12 3 15 INVX1
* cell instance $5 r0 *1 10.1,0
X$5 12 5 15 12 4 15 INVX1
* cell instance $6 r0 *1 11.9,0
X$6 12 6 15 12 5 15 INVX1
* cell instance $7 r0 *1 13.7,0
X$7 12 7 15 12 6 15 INVX1
* cell instance $8 r0 *1 15.5,0
X$8 12 8 15 12 7 15 INVX1
* cell instance $9 r0 *1 17.3,0
X$9 12 9 15 12 8 15 INVX1
* cell instance $10 r0 *1 19.1,0
X$10 12 10 15 12 9 15 INVX1
* cell instance $11 r0 *1 20.9,0
X$11 12 11 15 12 10 15 INVX1
* cell instance $12 r0 *1 24.7,0
X$12 12 13 15 12 11 15 INVX1
.ENDS RINGO

* cell INVX1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin IN
* pin SUBSTRATE
.SUBCKT INVX1 1 2 3 4 5 6
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 IN
* net 6 SUBSTRATE
* device instance $1 r0 *1 0.85,5.8 PMOS
M$1 1 5 2 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $2 r0 *1 0.85,2.135 NMOS
M$2 3 5 2 6 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
.ENDS INVX1

* cell ND2X1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin B
* pin A
* pin SUBSTRATE
.SUBCKT ND2X1 1 2 3 4 5 6 7
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 B
* net 6 A
* net 7 SUBSTRATE
* device instance $1 r0 *1 0.85,5.8 PMOS
M$1 2 6 1 4 PMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 r0 *1 1.55,5.8 PMOS
M$2 1 5 2 4 PMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 r0 *1 0.85,2.135 NMOS
M$3 3 6 8 7 NMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U PD=1.4U
* device instance $4 r0 *1 1.55,2.135 NMOS
M$4 8 5 2 7 NMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
.ENDS ND2X1
