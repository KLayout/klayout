magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 504 216 540
rect 324 504 468 540
rect 0 468 504 504
rect 0 396 540 468
rect 0 0 108 396
rect 216 0 324 396
rect 432 0 540 396
<< properties >>
string FIXED_BBOX 0 -216 648 756
<< end >>
