magic
tech scmos
timestamp 1534325869
<< silk >>
rect 0 8 12 12
<< end >>
