VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.002 ;

USEMINSPACING OBS OFF ;

END LIBRARY

LAYER overlap
	TYPE OVERLAP ;
END overlap

LAYER contact
	TYPE CUT ;
END contact

END LIBRARY

LAYER metal1
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
END metal1

LAYER via1
	TYPE CUT ;
END via1

LAYER metal2
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
END metal2

LAYER via2
	TYPE CUT ;
END via2

LAYER metal3
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
END metal3

LAYER via3
	TYPE CUT ;
END via3

LAYER metal4
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
END metal4

END LIBRARY
LAYER via4
	TYPE CUT ;
END via4

LAYER metal5
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
END metal5

END LIBRARY
