* netlist

* cell TOP1
.SUBCKT TOP1
.ENDS TOP1
