magic
tech scmos
timestamp 1540544905
<< polysilicon >>
rect 147 161 152 168
rect 147 130 152 137
<< metal1 >>
rect 90 178 100 200
rect 200 178 210 200
rect 90 168 145 178
rect 155 168 210 178
rect 90 120 145 130
rect 155 120 210 130
rect 90 100 100 120
rect 200 100 210 120
<< rnfet >>
rect 147 144 152 148
<< rpfet >>
rect 147 150 152 154
<< rpoly >>
rect 147 148 152 150
<< polycontact >>
rect 145 168 155 178
rect 145 120 155 130
<< polyndiff >>
rect 147 137 152 144
<< polypdiff >>
rect 147 154 152 161
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_k  L500_CHAR_k_0
timestamp 1534322894
transform 1 0 145 0 1 260
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 225 0 1 140
box 0 0 12 18
use Library/magic/L500_CHAR_w  L500_CHAR_w_0
timestamp 1534324213
transform 1 0 244 0 1 151
box 0 0 16 18
use Library/magic/L500_CHAR_5  L500_CHAR_5_0
timestamp 1534324893
transform 1 0 264 0 1 151
box 0 0 12 18
use Library/magic/L500_CHAR_slash  L500_CHAR_slash_0
timestamp 1534532558
transform 1 0 280 0 1 151
box 0 0 8 18
use Library/magic/L500_CHAR_l  L500_CHAR_l_0
timestamp 1534225390
transform 1 0 244 0 1 129
box 0 0 12 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_1
timestamp 1534324708
transform 1 0 260 0 1 129
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 145 0 1 20
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
