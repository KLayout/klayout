magic
tech scmos
timestamp 1534327094
<< silk >>
rect 0 8 4 18
rect 0 0 4 4
<< end >>
