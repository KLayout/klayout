UNITS
  DATABASE MICRONS 1000 ;
END UNITS
END LIBRARY
