VERSION 5.8 ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.1 ;
  PITCH 0.1 ;
END M1

LAYER overlap
  TYPE OVERLAP ;
END overlap
