magic
tech scmos
timestamp 1534325357
<< silk >>
rect 4 17 12 18
rect 2 16 12 17
rect 1 14 12 16
rect 0 13 5 14
rect 0 10 4 13
rect 8 10 12 14
rect 0 6 12 10
rect 0 0 4 6
rect 8 0 12 6
<< end >>
