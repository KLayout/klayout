VERSION 5.4 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
NOWIREEXTENSIONATPIN OFF ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER M1
    TYPE ROUTING ;
END M1

LAYER VIA1
    TYPE CUT ;
END VIA1

LAYER M2
    TYPE ROUTING ;
END M2

END LIBRARY
