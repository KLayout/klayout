UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

LAYER M1
  TYPE ROUTING ;
  WIDTH 0.002 ;
END M1

