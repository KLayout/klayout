magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 648 108 756
rect 432 648 540 756
rect 0 540 216 648
rect 324 540 540 648
rect 0 432 540 540
rect 0 0 108 432
rect 216 324 324 432
rect 432 0 540 432
<< properties >>
string FIXED_BBOX 0 -216 648 756
<< end >>
