magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 0 216 216
rect 108 -108 216 0
<< properties >>
string FIXED_BBOX 0 -216 324 756
<< end >>
