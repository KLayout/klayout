magic
timestamp 1575832387
<< checkpaint >>
rect -1 -3 12 18
<< l5d0 >>
rect 4 -3 7 18
rect 4 -3 7 18
<< l1001d0 >>
rect 8 1 11 15
rect 1 1 4 15
<< l2d0 >>
rect 0 0 11 15
rect 0 0 11 15
<< l1000d0 >>
rect 1 7 3 8
rect 8 7 10 8
rect 1 1 3 3
rect 8 1 10 3
rect 8 12 10 14
rect 1 12 3 14
<< l3d0 >>
rect -1 -1 12 16
<< end >>
