magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 720 252 756
rect 0 684 288 720
rect 0 612 324 684
rect 0 504 108 612
rect 216 504 324 612
rect 0 432 324 504
rect 0 396 288 432
rect 0 360 252 396
rect 0 252 216 360
rect 0 216 252 252
rect 0 180 288 216
rect 0 108 324 180
rect 0 0 108 108
rect 216 0 324 108
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
