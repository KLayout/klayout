magic
tech scmos
timestamp 1541639606
<< metal1 >>
rect 100 205 101 206
rect 199 205 200 206
rect 100 204 102 205
rect 198 204 200 205
rect 100 203 103 204
rect 197 203 200 204
rect 100 202 104 203
rect 196 202 200 203
rect 100 201 105 202
rect 195 201 200 202
rect 100 200 106 201
rect 194 200 200 201
rect 95 199 107 200
rect 193 199 205 200
rect 96 198 108 199
rect 192 198 204 199
rect 97 197 109 198
rect 191 197 203 198
rect 98 196 110 197
rect 190 196 202 197
rect 99 195 111 196
rect 189 195 201 196
rect 100 194 112 195
rect 188 194 200 195
rect 101 193 113 194
rect 187 193 199 194
rect 102 192 114 193
rect 186 192 198 193
rect 103 191 115 192
rect 185 191 197 192
rect 104 190 116 191
rect 184 190 196 191
rect 105 189 117 190
rect 183 189 195 190
rect 106 188 118 189
rect 182 188 194 189
rect 107 187 119 188
rect 181 187 193 188
rect 108 186 120 187
rect 180 186 192 187
rect 109 185 121 186
rect 179 185 191 186
rect 110 184 122 185
rect 178 184 190 185
rect 111 183 123 184
rect 177 183 189 184
rect 112 182 124 183
rect 176 182 188 183
rect 113 181 125 182
rect 175 181 187 182
rect 114 180 126 181
rect 174 180 186 181
rect 115 179 127 180
rect 173 179 185 180
rect 116 178 128 179
rect 172 178 184 179
rect 117 177 129 178
rect 171 177 183 178
rect 118 176 130 177
rect 170 176 182 177
rect 119 175 131 176
rect 169 175 181 176
rect 120 174 132 175
rect 168 174 180 175
rect 121 173 133 174
rect 167 173 179 174
rect 122 172 134 173
rect 166 172 178 173
rect 123 171 135 172
rect 165 171 177 172
rect 124 170 136 171
rect 164 170 176 171
rect 125 169 137 170
rect 163 169 175 170
rect 126 168 138 169
rect 162 168 174 169
rect 127 167 139 168
rect 161 167 173 168
rect 128 166 140 167
rect 160 166 172 167
rect 129 165 141 166
rect 159 165 171 166
rect 130 164 142 165
rect 158 164 170 165
rect 131 163 143 164
rect 157 163 169 164
rect 132 162 144 163
rect 156 162 168 163
rect 133 161 145 162
rect 155 161 167 162
rect 134 160 146 161
rect 154 160 166 161
rect 135 159 147 160
rect 153 159 165 160
rect 136 158 148 159
rect 137 157 148 158
rect 138 156 148 157
rect 139 155 148 156
rect 140 154 148 155
rect 141 153 148 154
rect 152 158 164 159
rect 152 157 163 158
rect 152 156 162 157
rect 152 155 161 156
rect 152 154 160 155
rect 152 153 159 154
rect 142 152 158 153
rect 143 151 148 152
rect 144 150 148 151
rect 145 149 148 150
rect 146 148 148 149
rect 152 151 157 152
rect 152 150 156 151
rect 152 149 155 150
rect 152 148 154 149
rect 147 147 153 148
<< metal2 >>
rect 147 152 153 153
rect 146 151 148 152
rect 145 150 148 151
rect 144 149 148 150
rect 143 148 148 149
rect 152 151 154 152
rect 152 150 155 151
rect 152 149 156 150
rect 152 148 157 149
rect 142 147 158 148
rect 141 146 148 147
rect 140 145 148 146
rect 139 144 148 145
rect 138 143 148 144
rect 137 142 148 143
rect 136 141 148 142
rect 152 146 159 147
rect 152 145 160 146
rect 152 144 161 145
rect 152 143 162 144
rect 152 142 163 143
rect 152 141 164 142
rect 135 140 147 141
rect 153 140 165 141
rect 134 139 146 140
rect 154 139 166 140
rect 133 138 145 139
rect 155 138 167 139
rect 132 137 144 138
rect 156 137 168 138
rect 131 136 143 137
rect 157 136 169 137
rect 130 135 142 136
rect 158 135 170 136
rect 129 134 141 135
rect 159 134 171 135
rect 128 133 140 134
rect 160 133 172 134
rect 127 132 139 133
rect 161 132 173 133
rect 126 131 138 132
rect 162 131 174 132
rect 125 130 137 131
rect 163 130 175 131
rect 124 129 136 130
rect 164 129 176 130
rect 123 128 135 129
rect 165 128 177 129
rect 122 127 134 128
rect 166 127 178 128
rect 121 126 133 127
rect 167 126 179 127
rect 120 125 132 126
rect 168 125 180 126
rect 119 124 131 125
rect 169 124 181 125
rect 118 123 130 124
rect 170 123 182 124
rect 117 122 129 123
rect 171 122 183 123
rect 116 121 128 122
rect 172 121 184 122
rect 115 120 127 121
rect 173 120 185 121
rect 114 119 126 120
rect 174 119 186 120
rect 113 118 125 119
rect 175 118 187 119
rect 112 117 124 118
rect 176 117 188 118
rect 111 116 123 117
rect 177 116 189 117
rect 110 115 122 116
rect 178 115 190 116
rect 109 114 121 115
rect 179 114 191 115
rect 108 113 120 114
rect 180 113 192 114
rect 107 112 119 113
rect 181 112 193 113
rect 106 111 118 112
rect 182 111 194 112
rect 105 110 117 111
rect 183 110 195 111
rect 104 109 116 110
rect 184 109 196 110
rect 103 108 115 109
rect 185 108 197 109
rect 102 107 114 108
rect 186 107 198 108
rect 101 106 113 107
rect 187 106 199 107
rect 100 105 112 106
rect 188 105 200 106
rect 99 104 111 105
rect 189 104 201 105
rect 98 103 110 104
rect 190 103 202 104
rect 97 102 109 103
rect 191 102 203 103
rect 96 101 108 102
rect 192 101 204 102
rect 95 100 107 101
rect 193 100 205 101
rect 100 99 106 100
rect 194 99 200 100
rect 100 98 105 99
rect 195 98 200 99
rect 100 97 104 98
rect 196 97 200 98
rect 100 96 103 97
rect 197 96 200 97
rect 100 95 102 96
rect 198 95 200 96
rect 100 94 101 95
rect 199 94 200 95
<< m2contact >>
rect 148 148 152 152
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_1
timestamp 1537343441
transform 1 0 0 0 1 200
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_3
timestamp 1537343441
transform 1 0 200 0 1 200
box 0 0 100 100
use Library/magic/L500_CHAR_m  L500_CHAR_m_2
timestamp 1534323034
transform 1 0 58 0 1 178
box 0 0 16 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_0
timestamp 1534326485
transform 1 0 78 0 1 178
box 0 0 12 18
use Library/magic/L500_CHAR_m  L500_CHAR_m_3
timestamp 1534323034
transform 1 0 209 0 1 178
box 0 0 16 18
use Library/magic/L500_CHAR_1  L500_CHAR_1_1
timestamp 1534326485
transform 1 0 229 0 1 178
box 0 0 12 18
use Library/magic/L500_CHAR_v  L500_CHAR_v_0
timestamp 1534326655
transform 1 0 172 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_i  L500_CHAR_i_0
timestamp 1534226087
transform 1 0 188 0 1 141
box 0 0 8 18
use Library/magic/L500_CHAR_a  L500_CHAR_a_0
timestamp 1534325357
transform 1 0 200 0 1 141
box 0 0 12 18
use Library/magic/L500_CHAR_m  L500_CHAR_m_1
timestamp 1534323034
transform 1 0 58 0 1 104
box 0 0 16 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_1
timestamp 1534324708
transform 1 0 79 0 1 104
box 0 0 12 18
use Library/magic/L500_CHAR_m  L500_CHAR_m_0
timestamp 1534323034
transform 1 0 209 0 1 104
box 0 0 16 18
use Library/magic/L500_CHAR_2  L500_CHAR_2_0
timestamp 1534324708
transform 1 0 229 0 1 104
box 0 0 12 18
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_0
timestamp 1537343441
transform 1 0 0 0 1 0
box 0 0 100 100
use Library/magic/L500_TPAD_blank  L500_TPAD_blank_2
timestamp 1537343441
transform 1 0 200 0 1 0
box 0 0 100 100
<< end >>
