magic
tech scmos
timestamp 1534324947
<< silk >>
rect 1 16 12 18
rect 0 15 12 16
rect 0 12 4 15
rect 0 11 10 12
rect 0 10 11 11
rect 0 8 12 10
rect 0 4 4 8
rect 8 4 12 8
rect 0 2 12 4
rect 1 1 11 2
rect 2 0 10 1
<< end >>
