magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 504 108 756
rect 216 504 324 756
rect 0 432 324 504
rect 36 360 288 432
rect 72 288 252 360
rect 108 0 216 288
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
