magic
tech gf180mcuD
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 144 108 540
rect 216 144 324 540
rect 432 144 540 540
rect 0 72 540 144
rect 36 36 540 72
rect 72 0 216 36
rect 324 0 540 36
<< properties >>
string FIXED_BBOX 0 -216 648 756
<< end >>
