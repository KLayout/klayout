magic
tech scmos
timestamp 1534326655
<< silk >>
rect 0 13 3 18
rect 9 13 12 18
rect 0 10 4 13
rect 1 7 4 10
rect 8 10 12 13
rect 8 7 11 10
rect 1 4 11 7
rect 2 3 10 4
rect 3 1 9 3
rect 4 0 8 1
<< end >>
