magic
tech scmos
timestamp 1538544897
use Library/magic/L500_CHAR_v  L500_CHAR_v_0
timestamp 1534326655
transform 1 0 0 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_0
timestamp 1534321738
transform 1 0 16 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_d  L500_CHAR_d_1
timestamp 1534321738
transform 1 0 32 0 1 0
box 0 0 12 18
use Library/magic/L500_CHAR_mark  L500_CHAR_mark_0
timestamp 1534327094
transform 1 0 48 0 1 0
box 0 0 4 18
<< end >>
