magic
tech gf180mcuD
timestamp 1654634570
<< properties >>
string FIXED_BBOX 0 -43 86 151
<< end >>
