* RINGO netlist after simplification

* cell RINGO
* pin OUT
* pin ENABLE
* pin VDD
* pin FB
* pin BULK,VSS
.SUBCKT RINGO 11 13 14 15 16
* net 11 OUT
* net 13 ENABLE
* net 14 VDD
* net 15 FB
* net 16 BULK,VSS
* device instance $1 2.65,5.8 LVPMOS
M$1 1 13 14 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 3.35,5.8 LVPMOS
M$2 14 15 1 14 LVPMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 5.05,5.8 LVPMOS
M$3 14 1 2 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $4 6.85,5.8 LVPMOS
M$4 14 2 3 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $5 8.65,5.8 LVPMOS
M$5 14 3 4 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $6 10.45,5.8 LVPMOS
M$6 14 4 5 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $7 12.25,5.8 LVPMOS
M$7 14 5 6 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $8 14.05,5.8 LVPMOS
M$8 14 6 7 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $9 15.85,5.8 LVPMOS
M$9 14 7 8 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $10 17.65,5.8 LVPMOS
M$10 14 8 9 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $11 19.45,5.8 LVPMOS
M$11 14 9 10 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $12 21.25,5.8 LVPMOS
M$12 14 10 15 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $13 23.05,5.8 LVPMOS
M$13 14 15 11 14 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $14 2.65,2.135 LVNMOS
M$14 16 13 12 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U
+ PD=1.4U
* device instance $15 3.35,2.135 LVNMOS
M$15 12 15 1 16 LVNMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
* device instance $16 5.05,2.135 LVNMOS
M$16 16 1 2 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $17 6.85,2.135 LVNMOS
M$17 16 2 3 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $18 8.65,2.135 LVNMOS
M$18 16 3 4 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $19 10.45,2.135 LVNMOS
M$19 16 4 5 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $20 12.25,2.135 LVNMOS
M$20 16 5 6 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $21 14.05,2.135 LVNMOS
M$21 16 6 7 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $22 15.85,2.135 LVNMOS
M$22 16 7 8 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $23 17.65,2.135 LVNMOS
M$23 16 8 9 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
* device instance $24 19.45,2.135 LVNMOS
M$24 16 9 10 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
* device instance $25 21.25,2.135 LVNMOS
M$25 16 10 15 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
* device instance $26 23.05,2.135 LVNMOS
M$26 16 15 11 16 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U
+ PD=2.75U
.ENDS RINGO
