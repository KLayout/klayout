magic
timestamp 1575832387
<< checkpaint >>
rect -1 -3 12 12
<< l5d0 >>
rect 4 -3 7 12
<< l1001d0 >>
rect 8 1 11 9
rect 1 1 4 9
<< l2d0 >>
rect 0 0 11 10
<< l1000d0 >>
rect 1 7 3 8
rect 1 1 3 3
rect 8 1 10 3
rect 8 7 10 8
<< l4d0 >>
rect -1 -1 12 10
<< end >>
