VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
 
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;
 
LAYER METAL_1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
    WIDTH 0.6 ;
END METAL_1

LAYER VIA_1
  TYPE CUT ;
END VIA_1

LAYER METAL_2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
    WIDTH 0.6 ;
END METAL_2 

END LIBRARY

