MACRO macro1
    CLASS CORE ;
    FOREIGN foreign1  0.5 -0.2 W ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.384 BY 0.480 ;
    PIN Z
        PORT
        LAYER M1 ;
        RECT  0.306 0.357 0.318 0.403 ;
        RECT  0.318 0.115 0.352 0.403 ;
        VIA  0.336 0.167 square ;
        VIA  0.336 0.351 square ;
        END
    END Z
END macro1

MACRO macro2
    CLASS CORE ;
    FOREIGN foreign2  -0.15 0.25 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.384 BY 0.480 ;
    PIN Z
        PORT
        LAYER M1 ;
        RECT  0.306 0.357 0.318 0.403 ;
        RECT  0.318 0.115 0.352 0.403 ;
        VIA  0.336 0.167 square ;
        VIA  0.336 0.351 square ;
        END
    END Z
END macro2

MACRO macro3
    CLASS CORE ;
    FOREIGN macro3 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.384 BY 0.480 ;
    PIN Z
        PORT
        LAYER M1 ;
        RECT  0.306 0.357 0.318 0.403 ;
        RECT  0.318 0.115 0.352 0.403 ;
        VIA  0.336 0.167 square ;
        VIA  0.336 0.351 square ;
        END
    END Z
END macro3

