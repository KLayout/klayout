
* cell INVCHAIN
.SUBCKT INVCHAIN
X$1 9 7 8 6 9 5 1 5 3 2 13 14 INV3
X$2 8 11 9 10 8 11 2 12 2 12 5 4 13 14 INV2
X$3 14 13 11 12 4 4 10 10 INV
.ENDS INVCHAIN

* cell INV3
.SUBCKT INV3 1 2 3 4 5 6 7 8 9 10 11 12
X$1 12 11 3 10 8 6 1 5 INV
X$2 12 11 4 7 9 9 2 2 INV
X$3 12 11 2 9 7 7 4 4 INV
.ENDS INV3

* cell INV2
.SUBCKT INV2 1 2 3 4 5 6 7 8 9 10 11 12 13 14
X$1 14 13 3 11 9 7 1 5 INV
X$2 14 13 4 12 10 8 2 6 INV
.ENDS INV2

* cell INV
.SUBCKT INV 1 2 3 4 5 6 7 8
M$1 4 3 2 4 PMOS L=0.25U W=0.95U AS=0.79325P AD=0.26125P PS=3.57U PD=1.5U
M$2 2 7 5 2 PMOS L=0.25U W=0.95U AS=0.26125P AD=0.03325P PS=1.5U PD=1.97U
M$3 4 3 1 4 NMOS L=0.25U W=0.95U AS=0.79325P AD=0.26125P PS=3.57U PD=1.5U
M$4 1 8 6 1 NMOS L=0.25U W=0.95U AS=0.26125P AD=0.03325P PS=1.5U PD=1.97U
.ENDS INV

