* VDIV netlist after simplification

* cell TOP
* pin OUT
* pin GND
* pin IN
* pin VDD
.SUBCKT TOP 1 2 3 5
* net 1 OUT
* net 2 GND
* net 3 IN
* net 5 VDD
* device instance $1 1.025,0.335 RES
R$1 4 1 7650
* device instance $2 2.85,0.335 RES
R$2 2 1 10320
* device instance $4 1.765,7.485 HVPMOS
M$4 4 3 5 5 MHVPMOS L=0.25U W=1.5U AS=0.63P AD=0.63P PS=3.84U PD=3.84U
.ENDS TOP
