
* cell INVCHAIN
.SUBCKT INVCHAIN
X$1 1 2 3 4 4 5 5 6 INV3
X$2 1 2 6 7 7 8 INV2
X$3 1 2 8 9 INV
.ENDS INVCHAIN

* cell INV3
.SUBCKT INV3 1 2 3 4 5 6 7 8 
X$1 1 2 3 4 INV
X$2 1 2 5 6 INV
X$3 1 2 7 8 INV
.ENDS INV3

* cell INV2
.SUBCKT INV2 1 2 3 4 5 6 
X$1 1 2 3 4 INV
X$2 1 2 5 6 INV
.ENDS INV2

* cell INV
.SUBCKT INV 1 2 3 4 
M$1 1 3 4 1 PMOS L=0.25U W=0.95U
M$3 2 3 4 2 NMOS L=0.25U W=0.95U
.ENDS INV

