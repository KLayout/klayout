* Extracted by KLayout

.SUBCKT TOP
X$1 \$2 \$5 \$4 E \$1 MIDDLE
.ENDS TOP

.SUBCKT MIDDLE B \$I4 \$I3 \$I2 \$I1
X$1 \$I1 B \$I3 \$I4 \$I2 F CHILD
.ENDS MIDDLE

.SUBCKT CHILD A B C D \$8 \$9
.ENDS CHILD
