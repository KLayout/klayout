.subckt INVX1 1 2 3 4 5 6
  .include nreader14x.cir
.ends 

