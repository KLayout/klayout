VERSION 5.6 ;

UNITS
DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
VIA OR_DEFAULT STRING ;
END PROPERTYDEFINITIONS

LAYER metal1
TYPE ROUTING ;
END metal1

LAYER via1
TYPE CUT ;
END via1

LAYER metal2
TYPE ROUTING ;
END metal2

VIA via1_4 DEFAULT
LAYER via1 ;
RECT -0.035 -0.035 0.035 0.035 ;
LAYER metal1 ;
RECT -0.035 -0.07 0.035 0.07 ;
LAYER metal2 ;
RECT -0.035 -0.07 0.035 0.07 ;
PROPERTY OR_DEFAULT Y ;
END via1_4

END LIBRARY
