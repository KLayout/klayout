magic
tech scmos
timestamp 1533657739
<< silk >>
rect 426 546 427 547
rect 427 546 428 547
rect 426 545 427 546
rect 427 545 428 546
rect 424 544 425 545
rect 425 544 426 545
rect 426 544 427 545
rect 427 544 428 545
rect 428 544 429 545
rect 429 544 430 545
rect 430 544 431 545
rect 431 544 432 545
rect 424 543 425 544
rect 425 543 426 544
rect 426 543 427 544
rect 427 543 428 544
rect 428 543 429 544
rect 429 543 430 544
rect 430 543 431 544
rect 431 543 432 544
rect 420 542 421 543
rect 421 542 422 543
rect 422 542 423 543
rect 423 542 424 543
rect 424 542 425 543
rect 425 542 426 543
rect 426 542 427 543
rect 427 542 428 543
rect 428 542 429 543
rect 429 542 430 543
rect 430 542 431 543
rect 431 542 432 543
rect 420 541 421 542
rect 421 541 422 542
rect 422 541 423 542
rect 423 541 424 542
rect 424 541 425 542
rect 425 541 426 542
rect 426 541 427 542
rect 427 541 428 542
rect 428 541 429 542
rect 429 541 430 542
rect 430 541 431 542
rect 431 541 432 542
rect 418 540 419 541
rect 419 540 420 541
rect 420 540 421 541
rect 421 540 422 541
rect 422 540 423 541
rect 423 540 424 541
rect 424 540 425 541
rect 425 540 426 541
rect 426 540 427 541
rect 427 540 428 541
rect 428 540 429 541
rect 429 540 430 541
rect 430 540 431 541
rect 431 540 432 541
rect 432 540 433 541
rect 433 540 434 541
rect 418 539 419 540
rect 419 539 420 540
rect 420 539 421 540
rect 421 539 422 540
rect 422 539 423 540
rect 423 539 424 540
rect 424 539 425 540
rect 425 539 426 540
rect 426 539 427 540
rect 427 539 428 540
rect 428 539 429 540
rect 429 539 430 540
rect 430 539 431 540
rect 431 539 432 540
rect 432 539 433 540
rect 433 539 434 540
rect 418 538 419 539
rect 419 538 420 539
rect 420 538 421 539
rect 421 538 422 539
rect 422 538 423 539
rect 423 538 424 539
rect 424 538 425 539
rect 425 538 426 539
rect 426 538 427 539
rect 427 538 428 539
rect 428 538 429 539
rect 429 538 430 539
rect 430 538 431 539
rect 431 538 432 539
rect 432 538 433 539
rect 433 538 434 539
rect 434 538 435 539
rect 435 538 436 539
rect 418 537 419 538
rect 419 537 420 538
rect 420 537 421 538
rect 421 537 422 538
rect 422 537 423 538
rect 423 537 424 538
rect 424 537 425 538
rect 425 537 426 538
rect 426 537 427 538
rect 427 537 428 538
rect 428 537 429 538
rect 429 537 430 538
rect 430 537 431 538
rect 431 537 432 538
rect 432 537 433 538
rect 433 537 434 538
rect 434 537 435 538
rect 435 537 436 538
rect 414 536 415 537
rect 415 536 416 537
rect 416 536 417 537
rect 417 536 418 537
rect 418 536 419 537
rect 419 536 420 537
rect 420 536 421 537
rect 421 536 422 537
rect 422 536 423 537
rect 423 536 424 537
rect 424 536 425 537
rect 425 536 426 537
rect 426 536 427 537
rect 427 536 428 537
rect 428 536 429 537
rect 429 536 430 537
rect 430 536 431 537
rect 431 536 432 537
rect 432 536 433 537
rect 433 536 434 537
rect 434 536 435 537
rect 435 536 436 537
rect 414 535 415 536
rect 415 535 416 536
rect 416 535 417 536
rect 417 535 418 536
rect 418 535 419 536
rect 419 535 420 536
rect 420 535 421 536
rect 421 535 422 536
rect 422 535 423 536
rect 423 535 424 536
rect 424 535 425 536
rect 425 535 426 536
rect 426 535 427 536
rect 427 535 428 536
rect 428 535 429 536
rect 429 535 430 536
rect 430 535 431 536
rect 431 535 432 536
rect 432 535 433 536
rect 433 535 434 536
rect 434 535 435 536
rect 435 535 436 536
rect 414 534 415 535
rect 415 534 416 535
rect 416 534 417 535
rect 417 534 418 535
rect 418 534 419 535
rect 419 534 420 535
rect 420 534 421 535
rect 421 534 422 535
rect 422 534 423 535
rect 423 534 424 535
rect 424 534 425 535
rect 425 534 426 535
rect 426 534 427 535
rect 427 534 428 535
rect 428 534 429 535
rect 429 534 430 535
rect 430 534 431 535
rect 431 534 432 535
rect 432 534 433 535
rect 433 534 434 535
rect 434 534 435 535
rect 435 534 436 535
rect 412 533 413 534
rect 413 533 414 534
rect 414 533 415 534
rect 415 533 416 534
rect 416 533 417 534
rect 417 533 418 534
rect 418 533 419 534
rect 419 533 420 534
rect 420 533 421 534
rect 421 533 422 534
rect 422 533 423 534
rect 423 533 424 534
rect 424 533 425 534
rect 425 533 426 534
rect 426 533 427 534
rect 427 533 428 534
rect 428 533 429 534
rect 429 533 430 534
rect 430 533 431 534
rect 431 533 432 534
rect 432 533 433 534
rect 433 533 434 534
rect 434 533 435 534
rect 435 533 436 534
rect 436 533 437 534
rect 437 533 438 534
rect 412 532 413 533
rect 413 532 414 533
rect 414 532 415 533
rect 415 532 416 533
rect 416 532 417 533
rect 417 532 418 533
rect 418 532 419 533
rect 419 532 420 533
rect 420 532 421 533
rect 421 532 422 533
rect 422 532 423 533
rect 423 532 424 533
rect 424 532 425 533
rect 425 532 426 533
rect 426 532 427 533
rect 427 532 428 533
rect 428 532 429 533
rect 429 532 430 533
rect 430 532 431 533
rect 431 532 432 533
rect 432 532 433 533
rect 433 532 434 533
rect 434 532 435 533
rect 435 532 436 533
rect 436 532 437 533
rect 437 532 438 533
rect 412 531 413 532
rect 413 531 414 532
rect 414 531 415 532
rect 415 531 416 532
rect 416 531 417 532
rect 417 531 418 532
rect 418 531 419 532
rect 419 531 420 532
rect 420 531 421 532
rect 421 531 422 532
rect 422 531 423 532
rect 423 531 424 532
rect 424 531 425 532
rect 425 531 426 532
rect 426 531 427 532
rect 427 531 428 532
rect 428 531 429 532
rect 429 531 430 532
rect 430 531 431 532
rect 431 531 432 532
rect 432 531 433 532
rect 433 531 434 532
rect 434 531 435 532
rect 435 531 436 532
rect 436 531 437 532
rect 437 531 438 532
rect 412 530 413 531
rect 413 530 414 531
rect 414 530 415 531
rect 415 530 416 531
rect 416 530 417 531
rect 417 530 418 531
rect 418 530 419 531
rect 419 530 420 531
rect 420 530 421 531
rect 421 530 422 531
rect 422 530 423 531
rect 423 530 424 531
rect 424 530 425 531
rect 425 530 426 531
rect 426 530 427 531
rect 427 530 428 531
rect 428 530 429 531
rect 429 530 430 531
rect 430 530 431 531
rect 431 530 432 531
rect 432 530 433 531
rect 433 530 434 531
rect 434 530 435 531
rect 435 530 436 531
rect 436 530 437 531
rect 437 530 438 531
rect 411 529 412 530
rect 412 529 413 530
rect 413 529 414 530
rect 414 529 415 530
rect 415 529 416 530
rect 416 529 417 530
rect 417 529 418 530
rect 418 529 419 530
rect 419 529 420 530
rect 420 529 421 530
rect 421 529 422 530
rect 422 529 423 530
rect 423 529 424 530
rect 424 529 425 530
rect 425 529 426 530
rect 426 529 427 530
rect 427 529 428 530
rect 428 529 429 530
rect 429 529 430 530
rect 430 529 431 530
rect 431 529 432 530
rect 432 529 433 530
rect 433 529 434 530
rect 434 529 435 530
rect 435 529 436 530
rect 436 529 437 530
rect 437 529 438 530
rect 411 528 412 529
rect 412 528 413 529
rect 413 528 414 529
rect 414 528 415 529
rect 415 528 416 529
rect 416 528 417 529
rect 417 528 418 529
rect 418 528 419 529
rect 419 528 420 529
rect 420 528 421 529
rect 421 528 422 529
rect 422 528 423 529
rect 423 528 424 529
rect 424 528 425 529
rect 425 528 426 529
rect 426 528 427 529
rect 427 528 428 529
rect 428 528 429 529
rect 429 528 430 529
rect 430 528 431 529
rect 431 528 432 529
rect 432 528 433 529
rect 433 528 434 529
rect 434 528 435 529
rect 435 528 436 529
rect 436 528 437 529
rect 437 528 438 529
rect 409 527 410 528
rect 410 527 411 528
rect 411 527 412 528
rect 412 527 413 528
rect 413 527 414 528
rect 414 527 415 528
rect 415 527 416 528
rect 416 527 417 528
rect 417 527 418 528
rect 418 527 419 528
rect 419 527 420 528
rect 420 527 421 528
rect 421 527 422 528
rect 422 527 423 528
rect 423 527 424 528
rect 424 527 425 528
rect 425 527 426 528
rect 426 527 427 528
rect 427 527 428 528
rect 428 527 429 528
rect 429 527 430 528
rect 430 527 431 528
rect 431 527 432 528
rect 432 527 433 528
rect 433 527 434 528
rect 434 527 435 528
rect 435 527 436 528
rect 436 527 437 528
rect 437 527 438 528
rect 438 527 439 528
rect 439 527 440 528
rect 409 526 410 527
rect 410 526 411 527
rect 411 526 412 527
rect 412 526 413 527
rect 413 526 414 527
rect 414 526 415 527
rect 415 526 416 527
rect 416 526 417 527
rect 417 526 418 527
rect 418 526 419 527
rect 419 526 420 527
rect 420 526 421 527
rect 421 526 422 527
rect 422 526 423 527
rect 423 526 424 527
rect 424 526 425 527
rect 425 526 426 527
rect 426 526 427 527
rect 427 526 428 527
rect 428 526 429 527
rect 429 526 430 527
rect 430 526 431 527
rect 431 526 432 527
rect 432 526 433 527
rect 433 526 434 527
rect 434 526 435 527
rect 435 526 436 527
rect 436 526 437 527
rect 437 526 438 527
rect 438 526 439 527
rect 439 526 440 527
rect 407 525 408 526
rect 408 525 409 526
rect 409 525 410 526
rect 410 525 411 526
rect 411 525 412 526
rect 412 525 413 526
rect 413 525 414 526
rect 414 525 415 526
rect 415 525 416 526
rect 416 525 417 526
rect 417 525 418 526
rect 418 525 419 526
rect 419 525 420 526
rect 420 525 421 526
rect 421 525 422 526
rect 422 525 423 526
rect 423 525 424 526
rect 424 525 425 526
rect 425 525 426 526
rect 426 525 427 526
rect 427 525 428 526
rect 428 525 429 526
rect 429 525 430 526
rect 430 525 431 526
rect 431 525 432 526
rect 432 525 433 526
rect 433 525 434 526
rect 434 525 435 526
rect 435 525 436 526
rect 436 525 437 526
rect 437 525 438 526
rect 438 525 439 526
rect 439 525 440 526
rect 407 524 408 525
rect 408 524 409 525
rect 409 524 410 525
rect 410 524 411 525
rect 411 524 412 525
rect 412 524 413 525
rect 413 524 414 525
rect 414 524 415 525
rect 415 524 416 525
rect 416 524 417 525
rect 417 524 418 525
rect 418 524 419 525
rect 419 524 420 525
rect 420 524 421 525
rect 421 524 422 525
rect 422 524 423 525
rect 423 524 424 525
rect 424 524 425 525
rect 425 524 426 525
rect 426 524 427 525
rect 427 524 428 525
rect 428 524 429 525
rect 429 524 430 525
rect 430 524 431 525
rect 431 524 432 525
rect 432 524 433 525
rect 433 524 434 525
rect 434 524 435 525
rect 435 524 436 525
rect 436 524 437 525
rect 437 524 438 525
rect 438 524 439 525
rect 439 524 440 525
rect 405 523 406 524
rect 406 523 407 524
rect 407 523 408 524
rect 408 523 409 524
rect 409 523 410 524
rect 410 523 411 524
rect 411 523 412 524
rect 412 523 413 524
rect 413 523 414 524
rect 414 523 415 524
rect 415 523 416 524
rect 416 523 417 524
rect 417 523 418 524
rect 418 523 419 524
rect 419 523 420 524
rect 420 523 421 524
rect 421 523 422 524
rect 422 523 423 524
rect 423 523 424 524
rect 424 523 425 524
rect 425 523 426 524
rect 426 523 427 524
rect 427 523 428 524
rect 428 523 429 524
rect 429 523 430 524
rect 430 523 431 524
rect 431 523 432 524
rect 432 523 433 524
rect 433 523 434 524
rect 434 523 435 524
rect 435 523 436 524
rect 436 523 437 524
rect 437 523 438 524
rect 438 523 439 524
rect 439 523 440 524
rect 405 522 406 523
rect 406 522 407 523
rect 407 522 408 523
rect 408 522 409 523
rect 409 522 410 523
rect 410 522 411 523
rect 411 522 412 523
rect 412 522 413 523
rect 413 522 414 523
rect 414 522 415 523
rect 415 522 416 523
rect 416 522 417 523
rect 417 522 418 523
rect 418 522 419 523
rect 419 522 420 523
rect 420 522 421 523
rect 421 522 422 523
rect 422 522 423 523
rect 423 522 424 523
rect 424 522 425 523
rect 425 522 426 523
rect 426 522 427 523
rect 427 522 428 523
rect 428 522 429 523
rect 429 522 430 523
rect 430 522 431 523
rect 431 522 432 523
rect 432 522 433 523
rect 433 522 434 523
rect 434 522 435 523
rect 435 522 436 523
rect 436 522 437 523
rect 437 522 438 523
rect 438 522 439 523
rect 439 522 440 523
rect 403 521 404 522
rect 404 521 405 522
rect 405 521 406 522
rect 406 521 407 522
rect 407 521 408 522
rect 408 521 409 522
rect 409 521 410 522
rect 410 521 411 522
rect 411 521 412 522
rect 412 521 413 522
rect 413 521 414 522
rect 414 521 415 522
rect 415 521 416 522
rect 416 521 417 522
rect 417 521 418 522
rect 418 521 419 522
rect 419 521 420 522
rect 420 521 421 522
rect 421 521 422 522
rect 422 521 423 522
rect 423 521 424 522
rect 424 521 425 522
rect 425 521 426 522
rect 426 521 427 522
rect 427 521 428 522
rect 428 521 429 522
rect 429 521 430 522
rect 430 521 431 522
rect 431 521 432 522
rect 432 521 433 522
rect 433 521 434 522
rect 434 521 435 522
rect 435 521 436 522
rect 436 521 437 522
rect 437 521 438 522
rect 438 521 439 522
rect 439 521 440 522
rect 440 521 441 522
rect 441 521 442 522
rect 403 520 404 521
rect 404 520 405 521
rect 405 520 406 521
rect 406 520 407 521
rect 407 520 408 521
rect 408 520 409 521
rect 409 520 410 521
rect 410 520 411 521
rect 411 520 412 521
rect 412 520 413 521
rect 413 520 414 521
rect 414 520 415 521
rect 415 520 416 521
rect 416 520 417 521
rect 417 520 418 521
rect 418 520 419 521
rect 419 520 420 521
rect 420 520 421 521
rect 421 520 422 521
rect 422 520 423 521
rect 423 520 424 521
rect 424 520 425 521
rect 425 520 426 521
rect 426 520 427 521
rect 427 520 428 521
rect 428 520 429 521
rect 429 520 430 521
rect 430 520 431 521
rect 431 520 432 521
rect 432 520 433 521
rect 433 520 434 521
rect 434 520 435 521
rect 435 520 436 521
rect 436 520 437 521
rect 437 520 438 521
rect 438 520 439 521
rect 439 520 440 521
rect 440 520 441 521
rect 441 520 442 521
rect 401 519 402 520
rect 402 519 403 520
rect 403 519 404 520
rect 404 519 405 520
rect 405 519 406 520
rect 406 519 407 520
rect 407 519 408 520
rect 408 519 409 520
rect 409 519 410 520
rect 410 519 411 520
rect 411 519 412 520
rect 412 519 413 520
rect 413 519 414 520
rect 414 519 415 520
rect 415 519 416 520
rect 416 519 417 520
rect 417 519 418 520
rect 418 519 419 520
rect 419 519 420 520
rect 420 519 421 520
rect 421 519 422 520
rect 422 519 423 520
rect 423 519 424 520
rect 424 519 425 520
rect 425 519 426 520
rect 426 519 427 520
rect 427 519 428 520
rect 428 519 429 520
rect 429 519 430 520
rect 430 519 431 520
rect 431 519 432 520
rect 432 519 433 520
rect 433 519 434 520
rect 434 519 435 520
rect 435 519 436 520
rect 436 519 437 520
rect 437 519 438 520
rect 438 519 439 520
rect 439 519 440 520
rect 440 519 441 520
rect 441 519 442 520
rect 401 518 402 519
rect 402 518 403 519
rect 403 518 404 519
rect 404 518 405 519
rect 405 518 406 519
rect 406 518 407 519
rect 407 518 408 519
rect 408 518 409 519
rect 409 518 410 519
rect 410 518 411 519
rect 411 518 412 519
rect 412 518 413 519
rect 413 518 414 519
rect 414 518 415 519
rect 415 518 416 519
rect 416 518 417 519
rect 417 518 418 519
rect 418 518 419 519
rect 419 518 420 519
rect 420 518 421 519
rect 421 518 422 519
rect 422 518 423 519
rect 423 518 424 519
rect 424 518 425 519
rect 425 518 426 519
rect 426 518 427 519
rect 427 518 428 519
rect 428 518 429 519
rect 429 518 430 519
rect 430 518 431 519
rect 431 518 432 519
rect 432 518 433 519
rect 433 518 434 519
rect 434 518 435 519
rect 435 518 436 519
rect 436 518 437 519
rect 437 518 438 519
rect 438 518 439 519
rect 439 518 440 519
rect 440 518 441 519
rect 441 518 442 519
rect 401 517 402 518
rect 402 517 403 518
rect 403 517 404 518
rect 404 517 405 518
rect 405 517 406 518
rect 406 517 407 518
rect 407 517 408 518
rect 408 517 409 518
rect 409 517 410 518
rect 410 517 411 518
rect 411 517 412 518
rect 412 517 413 518
rect 413 517 414 518
rect 414 517 415 518
rect 415 517 416 518
rect 416 517 417 518
rect 417 517 418 518
rect 418 517 419 518
rect 419 517 420 518
rect 420 517 421 518
rect 421 517 422 518
rect 422 517 423 518
rect 423 517 424 518
rect 424 517 425 518
rect 425 517 426 518
rect 426 517 427 518
rect 427 517 428 518
rect 428 517 429 518
rect 429 517 430 518
rect 430 517 431 518
rect 431 517 432 518
rect 432 517 433 518
rect 433 517 434 518
rect 434 517 435 518
rect 435 517 436 518
rect 436 517 437 518
rect 437 517 438 518
rect 438 517 439 518
rect 439 517 440 518
rect 440 517 441 518
rect 441 517 442 518
rect 401 516 402 517
rect 402 516 403 517
rect 403 516 404 517
rect 404 516 405 517
rect 405 516 406 517
rect 406 516 407 517
rect 407 516 408 517
rect 408 516 409 517
rect 409 516 410 517
rect 410 516 411 517
rect 411 516 412 517
rect 412 516 413 517
rect 413 516 414 517
rect 414 516 415 517
rect 415 516 416 517
rect 416 516 417 517
rect 417 516 418 517
rect 418 516 419 517
rect 419 516 420 517
rect 420 516 421 517
rect 421 516 422 517
rect 422 516 423 517
rect 423 516 424 517
rect 424 516 425 517
rect 425 516 426 517
rect 426 516 427 517
rect 427 516 428 517
rect 428 516 429 517
rect 429 516 430 517
rect 430 516 431 517
rect 431 516 432 517
rect 432 516 433 517
rect 433 516 434 517
rect 434 516 435 517
rect 435 516 436 517
rect 436 516 437 517
rect 437 516 438 517
rect 438 516 439 517
rect 439 516 440 517
rect 440 516 441 517
rect 441 516 442 517
rect 399 515 400 516
rect 400 515 401 516
rect 401 515 402 516
rect 402 515 403 516
rect 403 515 404 516
rect 404 515 405 516
rect 405 515 406 516
rect 406 515 407 516
rect 407 515 408 516
rect 408 515 409 516
rect 409 515 410 516
rect 410 515 411 516
rect 411 515 412 516
rect 412 515 413 516
rect 413 515 414 516
rect 414 515 415 516
rect 415 515 416 516
rect 416 515 417 516
rect 417 515 418 516
rect 418 515 419 516
rect 419 515 420 516
rect 420 515 421 516
rect 421 515 422 516
rect 422 515 423 516
rect 423 515 424 516
rect 424 515 425 516
rect 425 515 426 516
rect 426 515 427 516
rect 427 515 428 516
rect 428 515 429 516
rect 429 515 430 516
rect 430 515 431 516
rect 431 515 432 516
rect 432 515 433 516
rect 433 515 434 516
rect 434 515 435 516
rect 435 515 436 516
rect 436 515 437 516
rect 437 515 438 516
rect 438 515 439 516
rect 439 515 440 516
rect 440 515 441 516
rect 441 515 442 516
rect 399 514 400 515
rect 400 514 401 515
rect 401 514 402 515
rect 402 514 403 515
rect 403 514 404 515
rect 404 514 405 515
rect 405 514 406 515
rect 406 514 407 515
rect 407 514 408 515
rect 408 514 409 515
rect 409 514 410 515
rect 410 514 411 515
rect 411 514 412 515
rect 412 514 413 515
rect 413 514 414 515
rect 414 514 415 515
rect 415 514 416 515
rect 416 514 417 515
rect 417 514 418 515
rect 418 514 419 515
rect 419 514 420 515
rect 420 514 421 515
rect 421 514 422 515
rect 422 514 423 515
rect 423 514 424 515
rect 424 514 425 515
rect 425 514 426 515
rect 426 514 427 515
rect 427 514 428 515
rect 428 514 429 515
rect 429 514 430 515
rect 430 514 431 515
rect 431 514 432 515
rect 432 514 433 515
rect 433 514 434 515
rect 434 514 435 515
rect 435 514 436 515
rect 436 514 437 515
rect 437 514 438 515
rect 438 514 439 515
rect 439 514 440 515
rect 440 514 441 515
rect 441 514 442 515
rect 397 513 398 514
rect 398 513 399 514
rect 399 513 400 514
rect 400 513 401 514
rect 401 513 402 514
rect 402 513 403 514
rect 403 513 404 514
rect 404 513 405 514
rect 405 513 406 514
rect 406 513 407 514
rect 407 513 408 514
rect 408 513 409 514
rect 409 513 410 514
rect 410 513 411 514
rect 411 513 412 514
rect 412 513 413 514
rect 413 513 414 514
rect 414 513 415 514
rect 415 513 416 514
rect 416 513 417 514
rect 417 513 418 514
rect 418 513 419 514
rect 419 513 420 514
rect 420 513 421 514
rect 421 513 422 514
rect 422 513 423 514
rect 423 513 424 514
rect 424 513 425 514
rect 425 513 426 514
rect 426 513 427 514
rect 427 513 428 514
rect 428 513 429 514
rect 429 513 430 514
rect 430 513 431 514
rect 431 513 432 514
rect 432 513 433 514
rect 433 513 434 514
rect 434 513 435 514
rect 435 513 436 514
rect 436 513 437 514
rect 437 513 438 514
rect 438 513 439 514
rect 439 513 440 514
rect 440 513 441 514
rect 441 513 442 514
rect 397 512 398 513
rect 398 512 399 513
rect 399 512 400 513
rect 400 512 401 513
rect 401 512 402 513
rect 402 512 403 513
rect 403 512 404 513
rect 404 512 405 513
rect 405 512 406 513
rect 406 512 407 513
rect 407 512 408 513
rect 408 512 409 513
rect 409 512 410 513
rect 410 512 411 513
rect 411 512 412 513
rect 412 512 413 513
rect 413 512 414 513
rect 414 512 415 513
rect 415 512 416 513
rect 416 512 417 513
rect 417 512 418 513
rect 418 512 419 513
rect 419 512 420 513
rect 420 512 421 513
rect 421 512 422 513
rect 422 512 423 513
rect 423 512 424 513
rect 424 512 425 513
rect 425 512 426 513
rect 426 512 427 513
rect 427 512 428 513
rect 428 512 429 513
rect 429 512 430 513
rect 430 512 431 513
rect 431 512 432 513
rect 432 512 433 513
rect 433 512 434 513
rect 434 512 435 513
rect 435 512 436 513
rect 436 512 437 513
rect 437 512 438 513
rect 438 512 439 513
rect 439 512 440 513
rect 440 512 441 513
rect 441 512 442 513
rect 396 511 397 512
rect 397 511 398 512
rect 398 511 399 512
rect 399 511 400 512
rect 400 511 401 512
rect 401 511 402 512
rect 402 511 403 512
rect 403 511 404 512
rect 404 511 405 512
rect 405 511 406 512
rect 406 511 407 512
rect 407 511 408 512
rect 408 511 409 512
rect 409 511 410 512
rect 410 511 411 512
rect 411 511 412 512
rect 412 511 413 512
rect 413 511 414 512
rect 414 511 415 512
rect 415 511 416 512
rect 416 511 417 512
rect 417 511 418 512
rect 418 511 419 512
rect 419 511 420 512
rect 420 511 421 512
rect 421 511 422 512
rect 422 511 423 512
rect 423 511 424 512
rect 424 511 425 512
rect 425 511 426 512
rect 426 511 427 512
rect 427 511 428 512
rect 428 511 429 512
rect 429 511 430 512
rect 430 511 431 512
rect 431 511 432 512
rect 432 511 433 512
rect 433 511 434 512
rect 434 511 435 512
rect 435 511 436 512
rect 436 511 437 512
rect 437 511 438 512
rect 438 511 439 512
rect 439 511 440 512
rect 440 511 441 512
rect 441 511 442 512
rect 442 511 443 512
rect 396 510 397 511
rect 397 510 398 511
rect 398 510 399 511
rect 399 510 400 511
rect 400 510 401 511
rect 401 510 402 511
rect 402 510 403 511
rect 403 510 404 511
rect 404 510 405 511
rect 405 510 406 511
rect 406 510 407 511
rect 407 510 408 511
rect 408 510 409 511
rect 409 510 410 511
rect 410 510 411 511
rect 411 510 412 511
rect 412 510 413 511
rect 413 510 414 511
rect 414 510 415 511
rect 415 510 416 511
rect 416 510 417 511
rect 417 510 418 511
rect 418 510 419 511
rect 419 510 420 511
rect 420 510 421 511
rect 421 510 422 511
rect 422 510 423 511
rect 423 510 424 511
rect 424 510 425 511
rect 425 510 426 511
rect 426 510 427 511
rect 427 510 428 511
rect 428 510 429 511
rect 429 510 430 511
rect 430 510 431 511
rect 431 510 432 511
rect 432 510 433 511
rect 433 510 434 511
rect 434 510 435 511
rect 435 510 436 511
rect 436 510 437 511
rect 437 510 438 511
rect 438 510 439 511
rect 439 510 440 511
rect 440 510 441 511
rect 441 510 442 511
rect 442 510 443 511
rect 263 509 264 510
rect 264 509 265 510
rect 265 509 266 510
rect 266 509 267 510
rect 267 509 268 510
rect 268 509 269 510
rect 269 509 270 510
rect 270 509 271 510
rect 271 509 272 510
rect 272 509 273 510
rect 273 509 274 510
rect 274 509 275 510
rect 275 509 276 510
rect 276 509 277 510
rect 277 509 278 510
rect 278 509 279 510
rect 279 509 280 510
rect 280 509 281 510
rect 281 509 282 510
rect 283 509 284 510
rect 284 509 285 510
rect 285 509 286 510
rect 394 509 395 510
rect 395 509 396 510
rect 396 509 397 510
rect 397 509 398 510
rect 398 509 399 510
rect 399 509 400 510
rect 400 509 401 510
rect 401 509 402 510
rect 402 509 403 510
rect 403 509 404 510
rect 404 509 405 510
rect 405 509 406 510
rect 406 509 407 510
rect 407 509 408 510
rect 408 509 409 510
rect 409 509 410 510
rect 410 509 411 510
rect 411 509 412 510
rect 412 509 413 510
rect 413 509 414 510
rect 414 509 415 510
rect 415 509 416 510
rect 416 509 417 510
rect 417 509 418 510
rect 418 509 419 510
rect 419 509 420 510
rect 420 509 421 510
rect 421 509 422 510
rect 422 509 423 510
rect 423 509 424 510
rect 424 509 425 510
rect 425 509 426 510
rect 426 509 427 510
rect 427 509 428 510
rect 428 509 429 510
rect 429 509 430 510
rect 430 509 431 510
rect 431 509 432 510
rect 432 509 433 510
rect 433 509 434 510
rect 434 509 435 510
rect 435 509 436 510
rect 436 509 437 510
rect 437 509 438 510
rect 438 509 439 510
rect 439 509 440 510
rect 440 509 441 510
rect 441 509 442 510
rect 442 509 443 510
rect 263 508 264 509
rect 264 508 265 509
rect 265 508 266 509
rect 266 508 267 509
rect 267 508 268 509
rect 268 508 269 509
rect 269 508 270 509
rect 270 508 271 509
rect 271 508 272 509
rect 272 508 273 509
rect 273 508 274 509
rect 274 508 275 509
rect 275 508 276 509
rect 276 508 277 509
rect 277 508 278 509
rect 278 508 279 509
rect 279 508 280 509
rect 280 508 281 509
rect 281 508 282 509
rect 283 508 284 509
rect 284 508 285 509
rect 285 508 286 509
rect 394 508 395 509
rect 395 508 396 509
rect 396 508 397 509
rect 397 508 398 509
rect 398 508 399 509
rect 399 508 400 509
rect 400 508 401 509
rect 401 508 402 509
rect 402 508 403 509
rect 403 508 404 509
rect 404 508 405 509
rect 405 508 406 509
rect 406 508 407 509
rect 407 508 408 509
rect 408 508 409 509
rect 409 508 410 509
rect 410 508 411 509
rect 411 508 412 509
rect 412 508 413 509
rect 413 508 414 509
rect 414 508 415 509
rect 415 508 416 509
rect 416 508 417 509
rect 417 508 418 509
rect 418 508 419 509
rect 419 508 420 509
rect 420 508 421 509
rect 421 508 422 509
rect 422 508 423 509
rect 423 508 424 509
rect 424 508 425 509
rect 425 508 426 509
rect 426 508 427 509
rect 427 508 428 509
rect 428 508 429 509
rect 429 508 430 509
rect 430 508 431 509
rect 431 508 432 509
rect 432 508 433 509
rect 433 508 434 509
rect 434 508 435 509
rect 435 508 436 509
rect 436 508 437 509
rect 437 508 438 509
rect 438 508 439 509
rect 439 508 440 509
rect 440 508 441 509
rect 441 508 442 509
rect 253 507 254 508
rect 254 507 255 508
rect 255 507 256 508
rect 256 507 257 508
rect 257 507 258 508
rect 258 507 259 508
rect 259 507 260 508
rect 260 507 261 508
rect 261 507 262 508
rect 262 507 263 508
rect 263 507 264 508
rect 264 507 265 508
rect 265 507 266 508
rect 266 507 267 508
rect 267 507 268 508
rect 268 507 269 508
rect 269 507 270 508
rect 270 507 271 508
rect 271 507 272 508
rect 272 507 273 508
rect 273 507 274 508
rect 274 507 275 508
rect 275 507 276 508
rect 276 507 277 508
rect 277 507 278 508
rect 278 507 279 508
rect 279 507 280 508
rect 280 507 281 508
rect 281 507 282 508
rect 282 507 283 508
rect 283 507 284 508
rect 284 507 285 508
rect 285 507 286 508
rect 286 507 287 508
rect 287 507 288 508
rect 288 507 289 508
rect 289 507 290 508
rect 290 507 291 508
rect 291 507 292 508
rect 292 507 293 508
rect 293 507 294 508
rect 294 507 295 508
rect 295 507 296 508
rect 296 507 297 508
rect 297 507 298 508
rect 298 507 299 508
rect 299 507 300 508
rect 300 507 301 508
rect 392 507 393 508
rect 393 507 394 508
rect 394 507 395 508
rect 395 507 396 508
rect 396 507 397 508
rect 397 507 398 508
rect 398 507 399 508
rect 399 507 400 508
rect 400 507 401 508
rect 401 507 402 508
rect 402 507 403 508
rect 403 507 404 508
rect 404 507 405 508
rect 405 507 406 508
rect 406 507 407 508
rect 407 507 408 508
rect 408 507 409 508
rect 409 507 410 508
rect 410 507 411 508
rect 411 507 412 508
rect 412 507 413 508
rect 413 507 414 508
rect 414 507 415 508
rect 415 507 416 508
rect 416 507 417 508
rect 417 507 418 508
rect 418 507 419 508
rect 419 507 420 508
rect 420 507 421 508
rect 421 507 422 508
rect 422 507 423 508
rect 423 507 424 508
rect 424 507 425 508
rect 425 507 426 508
rect 426 507 427 508
rect 427 507 428 508
rect 428 507 429 508
rect 429 507 430 508
rect 430 507 431 508
rect 431 507 432 508
rect 432 507 433 508
rect 433 507 434 508
rect 434 507 435 508
rect 435 507 436 508
rect 436 507 437 508
rect 437 507 438 508
rect 438 507 439 508
rect 439 507 440 508
rect 440 507 441 508
rect 441 507 442 508
rect 442 507 443 508
rect 253 506 254 507
rect 254 506 255 507
rect 255 506 256 507
rect 256 506 257 507
rect 257 506 258 507
rect 258 506 259 507
rect 259 506 260 507
rect 260 506 261 507
rect 261 506 262 507
rect 262 506 263 507
rect 263 506 264 507
rect 264 506 265 507
rect 265 506 266 507
rect 266 506 267 507
rect 267 506 268 507
rect 268 506 269 507
rect 269 506 270 507
rect 270 506 271 507
rect 271 506 272 507
rect 272 506 273 507
rect 273 506 274 507
rect 274 506 275 507
rect 275 506 276 507
rect 276 506 277 507
rect 277 506 278 507
rect 278 506 279 507
rect 279 506 280 507
rect 280 506 281 507
rect 281 506 282 507
rect 282 506 283 507
rect 283 506 284 507
rect 284 506 285 507
rect 285 506 286 507
rect 286 506 287 507
rect 287 506 288 507
rect 288 506 289 507
rect 289 506 290 507
rect 290 506 291 507
rect 291 506 292 507
rect 292 506 293 507
rect 293 506 294 507
rect 294 506 295 507
rect 295 506 296 507
rect 296 506 297 507
rect 297 506 298 507
rect 298 506 299 507
rect 299 506 300 507
rect 300 506 301 507
rect 392 506 393 507
rect 393 506 394 507
rect 394 506 395 507
rect 395 506 396 507
rect 396 506 397 507
rect 397 506 398 507
rect 398 506 399 507
rect 399 506 400 507
rect 400 506 401 507
rect 401 506 402 507
rect 402 506 403 507
rect 403 506 404 507
rect 404 506 405 507
rect 405 506 406 507
rect 406 506 407 507
rect 407 506 408 507
rect 408 506 409 507
rect 409 506 410 507
rect 410 506 411 507
rect 411 506 412 507
rect 412 506 413 507
rect 413 506 414 507
rect 414 506 415 507
rect 415 506 416 507
rect 416 506 417 507
rect 417 506 418 507
rect 418 506 419 507
rect 419 506 420 507
rect 420 506 421 507
rect 421 506 422 507
rect 422 506 423 507
rect 423 506 424 507
rect 424 506 425 507
rect 425 506 426 507
rect 426 506 427 507
rect 427 506 428 507
rect 428 506 429 507
rect 429 506 430 507
rect 430 506 431 507
rect 431 506 432 507
rect 432 506 433 507
rect 433 506 434 507
rect 434 506 435 507
rect 435 506 436 507
rect 436 506 437 507
rect 437 506 438 507
rect 438 506 439 507
rect 439 506 440 507
rect 440 506 441 507
rect 441 506 442 507
rect 442 506 443 507
rect 248 505 249 506
rect 249 505 250 506
rect 250 505 251 506
rect 251 505 252 506
rect 252 505 253 506
rect 253 505 254 506
rect 254 505 255 506
rect 255 505 256 506
rect 256 505 257 506
rect 257 505 258 506
rect 258 505 259 506
rect 259 505 260 506
rect 260 505 261 506
rect 261 505 262 506
rect 262 505 263 506
rect 263 505 264 506
rect 264 505 265 506
rect 265 505 266 506
rect 266 505 267 506
rect 267 505 268 506
rect 268 505 269 506
rect 269 505 270 506
rect 270 505 271 506
rect 271 505 272 506
rect 272 505 273 506
rect 273 505 274 506
rect 274 505 275 506
rect 275 505 276 506
rect 276 505 277 506
rect 277 505 278 506
rect 278 505 279 506
rect 279 505 280 506
rect 280 505 281 506
rect 281 505 282 506
rect 282 505 283 506
rect 283 505 284 506
rect 284 505 285 506
rect 285 505 286 506
rect 286 505 287 506
rect 287 505 288 506
rect 288 505 289 506
rect 289 505 290 506
rect 290 505 291 506
rect 291 505 292 506
rect 292 505 293 506
rect 293 505 294 506
rect 294 505 295 506
rect 295 505 296 506
rect 296 505 297 506
rect 297 505 298 506
rect 298 505 299 506
rect 299 505 300 506
rect 300 505 301 506
rect 301 505 302 506
rect 302 505 303 506
rect 303 505 304 506
rect 304 505 305 506
rect 305 505 306 506
rect 306 505 307 506
rect 307 505 308 506
rect 308 505 309 506
rect 309 505 310 506
rect 390 505 391 506
rect 391 505 392 506
rect 392 505 393 506
rect 393 505 394 506
rect 394 505 395 506
rect 395 505 396 506
rect 396 505 397 506
rect 397 505 398 506
rect 398 505 399 506
rect 399 505 400 506
rect 400 505 401 506
rect 401 505 402 506
rect 402 505 403 506
rect 403 505 404 506
rect 404 505 405 506
rect 405 505 406 506
rect 406 505 407 506
rect 407 505 408 506
rect 408 505 409 506
rect 409 505 410 506
rect 410 505 411 506
rect 411 505 412 506
rect 412 505 413 506
rect 413 505 414 506
rect 414 505 415 506
rect 415 505 416 506
rect 416 505 417 506
rect 417 505 418 506
rect 418 505 419 506
rect 419 505 420 506
rect 420 505 421 506
rect 421 505 422 506
rect 422 505 423 506
rect 423 505 424 506
rect 424 505 425 506
rect 425 505 426 506
rect 426 505 427 506
rect 427 505 428 506
rect 428 505 429 506
rect 429 505 430 506
rect 430 505 431 506
rect 431 505 432 506
rect 432 505 433 506
rect 433 505 434 506
rect 434 505 435 506
rect 435 505 436 506
rect 436 505 437 506
rect 437 505 438 506
rect 438 505 439 506
rect 439 505 440 506
rect 440 505 441 506
rect 441 505 442 506
rect 442 505 443 506
rect 248 504 249 505
rect 249 504 250 505
rect 250 504 251 505
rect 251 504 252 505
rect 252 504 253 505
rect 253 504 254 505
rect 254 504 255 505
rect 255 504 256 505
rect 256 504 257 505
rect 257 504 258 505
rect 258 504 259 505
rect 259 504 260 505
rect 260 504 261 505
rect 261 504 262 505
rect 262 504 263 505
rect 263 504 264 505
rect 264 504 265 505
rect 265 504 266 505
rect 266 504 267 505
rect 267 504 268 505
rect 268 504 269 505
rect 269 504 270 505
rect 270 504 271 505
rect 271 504 272 505
rect 272 504 273 505
rect 273 504 274 505
rect 274 504 275 505
rect 275 504 276 505
rect 276 504 277 505
rect 277 504 278 505
rect 278 504 279 505
rect 279 504 280 505
rect 280 504 281 505
rect 281 504 282 505
rect 282 504 283 505
rect 283 504 284 505
rect 284 504 285 505
rect 285 504 286 505
rect 286 504 287 505
rect 287 504 288 505
rect 288 504 289 505
rect 289 504 290 505
rect 290 504 291 505
rect 291 504 292 505
rect 292 504 293 505
rect 293 504 294 505
rect 294 504 295 505
rect 295 504 296 505
rect 296 504 297 505
rect 297 504 298 505
rect 298 504 299 505
rect 299 504 300 505
rect 300 504 301 505
rect 301 504 302 505
rect 302 504 303 505
rect 303 504 304 505
rect 304 504 305 505
rect 305 504 306 505
rect 306 504 307 505
rect 307 504 308 505
rect 308 504 309 505
rect 309 504 310 505
rect 390 504 391 505
rect 391 504 392 505
rect 392 504 393 505
rect 393 504 394 505
rect 394 504 395 505
rect 395 504 396 505
rect 396 504 397 505
rect 397 504 398 505
rect 398 504 399 505
rect 399 504 400 505
rect 400 504 401 505
rect 401 504 402 505
rect 402 504 403 505
rect 403 504 404 505
rect 404 504 405 505
rect 405 504 406 505
rect 406 504 407 505
rect 407 504 408 505
rect 408 504 409 505
rect 409 504 410 505
rect 410 504 411 505
rect 411 504 412 505
rect 412 504 413 505
rect 413 504 414 505
rect 414 504 415 505
rect 415 504 416 505
rect 416 504 417 505
rect 417 504 418 505
rect 418 504 419 505
rect 419 504 420 505
rect 420 504 421 505
rect 421 504 422 505
rect 422 504 423 505
rect 423 504 424 505
rect 424 504 425 505
rect 425 504 426 505
rect 426 504 427 505
rect 427 504 428 505
rect 428 504 429 505
rect 429 504 430 505
rect 430 504 431 505
rect 431 504 432 505
rect 432 504 433 505
rect 433 504 434 505
rect 434 504 435 505
rect 435 504 436 505
rect 436 504 437 505
rect 437 504 438 505
rect 438 504 439 505
rect 439 504 440 505
rect 440 504 441 505
rect 441 504 442 505
rect 442 504 443 505
rect 244 503 245 504
rect 245 503 246 504
rect 246 503 247 504
rect 247 503 248 504
rect 248 503 249 504
rect 249 503 250 504
rect 250 503 251 504
rect 251 503 252 504
rect 252 503 253 504
rect 253 503 254 504
rect 254 503 255 504
rect 255 503 256 504
rect 256 503 257 504
rect 257 503 258 504
rect 258 503 259 504
rect 259 503 260 504
rect 260 503 261 504
rect 261 503 262 504
rect 262 503 263 504
rect 263 503 264 504
rect 264 503 265 504
rect 265 503 266 504
rect 266 503 267 504
rect 267 503 268 504
rect 268 503 269 504
rect 269 503 270 504
rect 270 503 271 504
rect 271 503 272 504
rect 272 503 273 504
rect 273 503 274 504
rect 274 503 275 504
rect 275 503 276 504
rect 276 503 277 504
rect 277 503 278 504
rect 278 503 279 504
rect 279 503 280 504
rect 280 503 281 504
rect 281 503 282 504
rect 282 503 283 504
rect 283 503 284 504
rect 284 503 285 504
rect 285 503 286 504
rect 286 503 287 504
rect 287 503 288 504
rect 288 503 289 504
rect 289 503 290 504
rect 290 503 291 504
rect 291 503 292 504
rect 292 503 293 504
rect 293 503 294 504
rect 294 503 295 504
rect 295 503 296 504
rect 296 503 297 504
rect 297 503 298 504
rect 298 503 299 504
rect 299 503 300 504
rect 300 503 301 504
rect 301 503 302 504
rect 302 503 303 504
rect 303 503 304 504
rect 304 503 305 504
rect 305 503 306 504
rect 306 503 307 504
rect 307 503 308 504
rect 308 503 309 504
rect 309 503 310 504
rect 310 503 311 504
rect 311 503 312 504
rect 312 503 313 504
rect 313 503 314 504
rect 314 503 315 504
rect 315 503 316 504
rect 317 503 318 504
rect 318 503 319 504
rect 319 503 320 504
rect 390 503 391 504
rect 391 503 392 504
rect 392 503 393 504
rect 393 503 394 504
rect 394 503 395 504
rect 395 503 396 504
rect 396 503 397 504
rect 397 503 398 504
rect 398 503 399 504
rect 399 503 400 504
rect 400 503 401 504
rect 401 503 402 504
rect 402 503 403 504
rect 403 503 404 504
rect 404 503 405 504
rect 405 503 406 504
rect 406 503 407 504
rect 407 503 408 504
rect 408 503 409 504
rect 409 503 410 504
rect 410 503 411 504
rect 411 503 412 504
rect 412 503 413 504
rect 413 503 414 504
rect 414 503 415 504
rect 415 503 416 504
rect 416 503 417 504
rect 417 503 418 504
rect 418 503 419 504
rect 419 503 420 504
rect 420 503 421 504
rect 421 503 422 504
rect 422 503 423 504
rect 423 503 424 504
rect 424 503 425 504
rect 425 503 426 504
rect 426 503 427 504
rect 427 503 428 504
rect 428 503 429 504
rect 429 503 430 504
rect 430 503 431 504
rect 431 503 432 504
rect 432 503 433 504
rect 433 503 434 504
rect 434 503 435 504
rect 435 503 436 504
rect 436 503 437 504
rect 437 503 438 504
rect 438 503 439 504
rect 439 503 440 504
rect 440 503 441 504
rect 441 503 442 504
rect 442 503 443 504
rect 244 502 245 503
rect 245 502 246 503
rect 246 502 247 503
rect 247 502 248 503
rect 248 502 249 503
rect 249 502 250 503
rect 250 502 251 503
rect 251 502 252 503
rect 252 502 253 503
rect 253 502 254 503
rect 254 502 255 503
rect 255 502 256 503
rect 256 502 257 503
rect 257 502 258 503
rect 258 502 259 503
rect 259 502 260 503
rect 260 502 261 503
rect 261 502 262 503
rect 262 502 263 503
rect 263 502 264 503
rect 264 502 265 503
rect 265 502 266 503
rect 266 502 267 503
rect 267 502 268 503
rect 268 502 269 503
rect 269 502 270 503
rect 270 502 271 503
rect 274 502 275 503
rect 275 502 276 503
rect 276 502 277 503
rect 278 502 279 503
rect 279 502 280 503
rect 281 502 282 503
rect 282 502 283 503
rect 283 502 284 503
rect 289 502 290 503
rect 290 502 291 503
rect 291 502 292 503
rect 292 502 293 503
rect 293 502 294 503
rect 294 502 295 503
rect 295 502 296 503
rect 296 502 297 503
rect 297 502 298 503
rect 298 502 299 503
rect 299 502 300 503
rect 300 502 301 503
rect 301 502 302 503
rect 302 502 303 503
rect 303 502 304 503
rect 304 502 305 503
rect 305 502 306 503
rect 306 502 307 503
rect 307 502 308 503
rect 308 502 309 503
rect 309 502 310 503
rect 310 502 311 503
rect 311 502 312 503
rect 312 502 313 503
rect 313 502 314 503
rect 314 502 315 503
rect 315 502 316 503
rect 317 502 318 503
rect 318 502 319 503
rect 319 502 320 503
rect 390 502 391 503
rect 391 502 392 503
rect 392 502 393 503
rect 393 502 394 503
rect 394 502 395 503
rect 395 502 396 503
rect 396 502 397 503
rect 397 502 398 503
rect 398 502 399 503
rect 399 502 400 503
rect 400 502 401 503
rect 401 502 402 503
rect 402 502 403 503
rect 403 502 404 503
rect 404 502 405 503
rect 405 502 406 503
rect 406 502 407 503
rect 407 502 408 503
rect 409 502 410 503
rect 410 502 411 503
rect 411 502 412 503
rect 412 502 413 503
rect 413 502 414 503
rect 414 502 415 503
rect 415 502 416 503
rect 416 502 417 503
rect 417 502 418 503
rect 418 502 419 503
rect 419 502 420 503
rect 420 502 421 503
rect 421 502 422 503
rect 422 502 423 503
rect 423 502 424 503
rect 424 502 425 503
rect 425 502 426 503
rect 426 502 427 503
rect 427 502 428 503
rect 428 502 429 503
rect 429 502 430 503
rect 430 502 431 503
rect 431 502 432 503
rect 432 502 433 503
rect 433 502 434 503
rect 434 502 435 503
rect 435 502 436 503
rect 436 502 437 503
rect 437 502 438 503
rect 438 502 439 503
rect 439 502 440 503
rect 440 502 441 503
rect 441 502 442 503
rect 240 501 241 502
rect 241 501 242 502
rect 242 501 243 502
rect 243 501 244 502
rect 244 501 245 502
rect 245 501 246 502
rect 246 501 247 502
rect 247 501 248 502
rect 248 501 249 502
rect 249 501 250 502
rect 250 501 251 502
rect 251 501 252 502
rect 252 501 253 502
rect 253 501 254 502
rect 254 501 255 502
rect 255 501 256 502
rect 256 501 257 502
rect 257 501 258 502
rect 258 501 259 502
rect 259 501 260 502
rect 260 501 261 502
rect 261 501 262 502
rect 262 501 263 502
rect 263 501 264 502
rect 264 501 265 502
rect 265 501 266 502
rect 266 501 267 502
rect 267 501 268 502
rect 268 501 269 502
rect 269 501 270 502
rect 270 501 271 502
rect 274 501 275 502
rect 275 501 276 502
rect 276 501 277 502
rect 278 501 279 502
rect 279 501 280 502
rect 281 501 282 502
rect 282 501 283 502
rect 283 501 284 502
rect 289 501 290 502
rect 290 501 291 502
rect 291 501 292 502
rect 292 501 293 502
rect 293 501 294 502
rect 294 501 295 502
rect 295 501 296 502
rect 296 501 297 502
rect 297 501 298 502
rect 298 501 299 502
rect 299 501 300 502
rect 300 501 301 502
rect 301 501 302 502
rect 302 501 303 502
rect 303 501 304 502
rect 304 501 305 502
rect 305 501 306 502
rect 306 501 307 502
rect 307 501 308 502
rect 308 501 309 502
rect 309 501 310 502
rect 310 501 311 502
rect 311 501 312 502
rect 312 501 313 502
rect 313 501 314 502
rect 314 501 315 502
rect 315 501 316 502
rect 316 501 317 502
rect 317 501 318 502
rect 318 501 319 502
rect 319 501 320 502
rect 320 501 321 502
rect 321 501 322 502
rect 322 501 323 502
rect 323 501 324 502
rect 324 501 325 502
rect 388 501 389 502
rect 389 501 390 502
rect 390 501 391 502
rect 391 501 392 502
rect 392 501 393 502
rect 393 501 394 502
rect 394 501 395 502
rect 395 501 396 502
rect 396 501 397 502
rect 397 501 398 502
rect 398 501 399 502
rect 399 501 400 502
rect 400 501 401 502
rect 401 501 402 502
rect 402 501 403 502
rect 403 501 404 502
rect 404 501 405 502
rect 405 501 406 502
rect 406 501 407 502
rect 407 501 408 502
rect 409 501 410 502
rect 410 501 411 502
rect 411 501 412 502
rect 412 501 413 502
rect 413 501 414 502
rect 414 501 415 502
rect 415 501 416 502
rect 416 501 417 502
rect 417 501 418 502
rect 418 501 419 502
rect 419 501 420 502
rect 420 501 421 502
rect 421 501 422 502
rect 422 501 423 502
rect 423 501 424 502
rect 424 501 425 502
rect 425 501 426 502
rect 426 501 427 502
rect 427 501 428 502
rect 428 501 429 502
rect 429 501 430 502
rect 430 501 431 502
rect 431 501 432 502
rect 432 501 433 502
rect 433 501 434 502
rect 434 501 435 502
rect 435 501 436 502
rect 436 501 437 502
rect 437 501 438 502
rect 438 501 439 502
rect 439 501 440 502
rect 440 501 441 502
rect 441 501 442 502
rect 442 501 443 502
rect 240 500 241 501
rect 241 500 242 501
rect 242 500 243 501
rect 243 500 244 501
rect 244 500 245 501
rect 245 500 246 501
rect 246 500 247 501
rect 247 500 248 501
rect 248 500 249 501
rect 249 500 250 501
rect 250 500 251 501
rect 251 500 252 501
rect 252 500 253 501
rect 253 500 254 501
rect 254 500 255 501
rect 255 500 256 501
rect 257 500 258 501
rect 258 500 259 501
rect 259 500 260 501
rect 304 500 305 501
rect 305 500 306 501
rect 306 500 307 501
rect 308 500 309 501
rect 309 500 310 501
rect 310 500 311 501
rect 311 500 312 501
rect 312 500 313 501
rect 313 500 314 501
rect 314 500 315 501
rect 315 500 316 501
rect 316 500 317 501
rect 317 500 318 501
rect 318 500 319 501
rect 319 500 320 501
rect 320 500 321 501
rect 321 500 322 501
rect 322 500 323 501
rect 323 500 324 501
rect 324 500 325 501
rect 388 500 389 501
rect 389 500 390 501
rect 390 500 391 501
rect 391 500 392 501
rect 392 500 393 501
rect 393 500 394 501
rect 394 500 395 501
rect 395 500 396 501
rect 396 500 397 501
rect 397 500 398 501
rect 398 500 399 501
rect 399 500 400 501
rect 400 500 401 501
rect 401 500 402 501
rect 402 500 403 501
rect 403 500 404 501
rect 404 500 405 501
rect 405 500 406 501
rect 411 500 412 501
rect 412 500 413 501
rect 413 500 414 501
rect 414 500 415 501
rect 415 500 416 501
rect 416 500 417 501
rect 417 500 418 501
rect 418 500 419 501
rect 419 500 420 501
rect 420 500 421 501
rect 421 500 422 501
rect 422 500 423 501
rect 423 500 424 501
rect 424 500 425 501
rect 425 500 426 501
rect 426 500 427 501
rect 427 500 428 501
rect 428 500 429 501
rect 429 500 430 501
rect 430 500 431 501
rect 431 500 432 501
rect 432 500 433 501
rect 433 500 434 501
rect 434 500 435 501
rect 435 500 436 501
rect 436 500 437 501
rect 437 500 438 501
rect 438 500 439 501
rect 439 500 440 501
rect 440 500 441 501
rect 441 500 442 501
rect 442 500 443 501
rect 236 499 237 500
rect 237 499 238 500
rect 238 499 239 500
rect 239 499 240 500
rect 240 499 241 500
rect 241 499 242 500
rect 242 499 243 500
rect 243 499 244 500
rect 244 499 245 500
rect 245 499 246 500
rect 246 499 247 500
rect 247 499 248 500
rect 248 499 249 500
rect 249 499 250 500
rect 250 499 251 500
rect 251 499 252 500
rect 252 499 253 500
rect 253 499 254 500
rect 254 499 255 500
rect 255 499 256 500
rect 257 499 258 500
rect 258 499 259 500
rect 259 499 260 500
rect 304 499 305 500
rect 305 499 306 500
rect 306 499 307 500
rect 308 499 309 500
rect 309 499 310 500
rect 310 499 311 500
rect 311 499 312 500
rect 312 499 313 500
rect 313 499 314 500
rect 314 499 315 500
rect 315 499 316 500
rect 316 499 317 500
rect 317 499 318 500
rect 318 499 319 500
rect 319 499 320 500
rect 320 499 321 500
rect 321 499 322 500
rect 322 499 323 500
rect 323 499 324 500
rect 324 499 325 500
rect 325 499 326 500
rect 326 499 327 500
rect 327 499 328 500
rect 328 499 329 500
rect 386 499 387 500
rect 387 499 388 500
rect 388 499 389 500
rect 389 499 390 500
rect 390 499 391 500
rect 391 499 392 500
rect 392 499 393 500
rect 393 499 394 500
rect 394 499 395 500
rect 395 499 396 500
rect 396 499 397 500
rect 397 499 398 500
rect 398 499 399 500
rect 399 499 400 500
rect 400 499 401 500
rect 401 499 402 500
rect 402 499 403 500
rect 403 499 404 500
rect 404 499 405 500
rect 405 499 406 500
rect 411 499 412 500
rect 412 499 413 500
rect 413 499 414 500
rect 414 499 415 500
rect 415 499 416 500
rect 416 499 417 500
rect 417 499 418 500
rect 418 499 419 500
rect 419 499 420 500
rect 420 499 421 500
rect 421 499 422 500
rect 422 499 423 500
rect 423 499 424 500
rect 424 499 425 500
rect 425 499 426 500
rect 426 499 427 500
rect 427 499 428 500
rect 428 499 429 500
rect 429 499 430 500
rect 430 499 431 500
rect 431 499 432 500
rect 432 499 433 500
rect 433 499 434 500
rect 434 499 435 500
rect 435 499 436 500
rect 436 499 437 500
rect 437 499 438 500
rect 438 499 439 500
rect 439 499 440 500
rect 440 499 441 500
rect 441 499 442 500
rect 442 499 443 500
rect 236 498 237 499
rect 237 498 238 499
rect 238 498 239 499
rect 239 498 240 499
rect 240 498 241 499
rect 241 498 242 499
rect 242 498 243 499
rect 243 498 244 499
rect 244 498 245 499
rect 245 498 246 499
rect 246 498 247 499
rect 247 498 248 499
rect 248 498 249 499
rect 311 498 312 499
rect 312 498 313 499
rect 313 498 314 499
rect 314 498 315 499
rect 315 498 316 499
rect 316 498 317 499
rect 317 498 318 499
rect 318 498 319 499
rect 319 498 320 499
rect 320 498 321 499
rect 321 498 322 499
rect 322 498 323 499
rect 323 498 324 499
rect 324 498 325 499
rect 325 498 326 499
rect 326 498 327 499
rect 327 498 328 499
rect 328 498 329 499
rect 386 498 387 499
rect 387 498 388 499
rect 388 498 389 499
rect 389 498 390 499
rect 390 498 391 499
rect 391 498 392 499
rect 392 498 393 499
rect 393 498 394 499
rect 394 498 395 499
rect 395 498 396 499
rect 396 498 397 499
rect 397 498 398 499
rect 398 498 399 499
rect 399 498 400 499
rect 400 498 401 499
rect 401 498 402 499
rect 411 498 412 499
rect 412 498 413 499
rect 413 498 414 499
rect 414 498 415 499
rect 415 498 416 499
rect 416 498 417 499
rect 417 498 418 499
rect 418 498 419 499
rect 419 498 420 499
rect 420 498 421 499
rect 421 498 422 499
rect 422 498 423 499
rect 423 498 424 499
rect 424 498 425 499
rect 425 498 426 499
rect 426 498 427 499
rect 427 498 428 499
rect 428 498 429 499
rect 429 498 430 499
rect 430 498 431 499
rect 431 498 432 499
rect 432 498 433 499
rect 433 498 434 499
rect 434 498 435 499
rect 435 498 436 499
rect 436 498 437 499
rect 437 498 438 499
rect 438 498 439 499
rect 439 498 440 499
rect 440 498 441 499
rect 441 498 442 499
rect 442 498 443 499
rect 235 497 236 498
rect 236 497 237 498
rect 237 497 238 498
rect 238 497 239 498
rect 239 497 240 498
rect 240 497 241 498
rect 241 497 242 498
rect 242 497 243 498
rect 243 497 244 498
rect 244 497 245 498
rect 245 497 246 498
rect 246 497 247 498
rect 247 497 248 498
rect 248 497 249 498
rect 311 497 312 498
rect 312 497 313 498
rect 313 497 314 498
rect 314 497 315 498
rect 315 497 316 498
rect 316 497 317 498
rect 317 497 318 498
rect 318 497 319 498
rect 319 497 320 498
rect 320 497 321 498
rect 321 497 322 498
rect 322 497 323 498
rect 323 497 324 498
rect 324 497 325 498
rect 325 497 326 498
rect 326 497 327 498
rect 327 497 328 498
rect 328 497 329 498
rect 329 497 330 498
rect 330 497 331 498
rect 384 497 385 498
rect 385 497 386 498
rect 386 497 387 498
rect 387 497 388 498
rect 388 497 389 498
rect 389 497 390 498
rect 390 497 391 498
rect 391 497 392 498
rect 392 497 393 498
rect 393 497 394 498
rect 394 497 395 498
rect 395 497 396 498
rect 396 497 397 498
rect 397 497 398 498
rect 398 497 399 498
rect 399 497 400 498
rect 400 497 401 498
rect 401 497 402 498
rect 411 497 412 498
rect 412 497 413 498
rect 413 497 414 498
rect 414 497 415 498
rect 415 497 416 498
rect 416 497 417 498
rect 417 497 418 498
rect 418 497 419 498
rect 419 497 420 498
rect 420 497 421 498
rect 421 497 422 498
rect 422 497 423 498
rect 423 497 424 498
rect 424 497 425 498
rect 425 497 426 498
rect 426 497 427 498
rect 427 497 428 498
rect 428 497 429 498
rect 429 497 430 498
rect 430 497 431 498
rect 431 497 432 498
rect 432 497 433 498
rect 433 497 434 498
rect 434 497 435 498
rect 435 497 436 498
rect 436 497 437 498
rect 437 497 438 498
rect 438 497 439 498
rect 439 497 440 498
rect 440 497 441 498
rect 441 497 442 498
rect 442 497 443 498
rect 235 496 236 497
rect 236 496 237 497
rect 237 496 238 497
rect 238 496 239 497
rect 239 496 240 497
rect 240 496 241 497
rect 241 496 242 497
rect 242 496 243 497
rect 317 496 318 497
rect 318 496 319 497
rect 319 496 320 497
rect 320 496 321 497
rect 321 496 322 497
rect 322 496 323 497
rect 323 496 324 497
rect 324 496 325 497
rect 325 496 326 497
rect 326 496 327 497
rect 327 496 328 497
rect 328 496 329 497
rect 329 496 330 497
rect 330 496 331 497
rect 384 496 385 497
rect 385 496 386 497
rect 386 496 387 497
rect 387 496 388 497
rect 388 496 389 497
rect 389 496 390 497
rect 390 496 391 497
rect 391 496 392 497
rect 392 496 393 497
rect 393 496 394 497
rect 394 496 395 497
rect 395 496 396 497
rect 396 496 397 497
rect 397 496 398 497
rect 398 496 399 497
rect 399 496 400 497
rect 412 496 413 497
rect 413 496 414 497
rect 414 496 415 497
rect 415 496 416 497
rect 416 496 417 497
rect 417 496 418 497
rect 418 496 419 497
rect 419 496 420 497
rect 420 496 421 497
rect 421 496 422 497
rect 422 496 423 497
rect 423 496 424 497
rect 424 496 425 497
rect 425 496 426 497
rect 426 496 427 497
rect 427 496 428 497
rect 428 496 429 497
rect 429 496 430 497
rect 430 496 431 497
rect 431 496 432 497
rect 432 496 433 497
rect 433 496 434 497
rect 434 496 435 497
rect 435 496 436 497
rect 436 496 437 497
rect 437 496 438 497
rect 438 496 439 497
rect 439 496 440 497
rect 440 496 441 497
rect 441 496 442 497
rect 442 496 443 497
rect 231 495 232 496
rect 232 495 233 496
rect 233 495 234 496
rect 234 495 235 496
rect 235 495 236 496
rect 236 495 237 496
rect 237 495 238 496
rect 238 495 239 496
rect 239 495 240 496
rect 240 495 241 496
rect 241 495 242 496
rect 242 495 243 496
rect 317 495 318 496
rect 318 495 319 496
rect 319 495 320 496
rect 320 495 321 496
rect 321 495 322 496
rect 322 495 323 496
rect 323 495 324 496
rect 324 495 325 496
rect 325 495 326 496
rect 326 495 327 496
rect 327 495 328 496
rect 328 495 329 496
rect 329 495 330 496
rect 330 495 331 496
rect 331 495 332 496
rect 332 495 333 496
rect 333 495 334 496
rect 334 495 335 496
rect 383 495 384 496
rect 384 495 385 496
rect 385 495 386 496
rect 386 495 387 496
rect 387 495 388 496
rect 388 495 389 496
rect 389 495 390 496
rect 390 495 391 496
rect 391 495 392 496
rect 392 495 393 496
rect 393 495 394 496
rect 394 495 395 496
rect 395 495 396 496
rect 396 495 397 496
rect 397 495 398 496
rect 398 495 399 496
rect 399 495 400 496
rect 412 495 413 496
rect 413 495 414 496
rect 414 495 415 496
rect 415 495 416 496
rect 416 495 417 496
rect 417 495 418 496
rect 418 495 419 496
rect 419 495 420 496
rect 420 495 421 496
rect 421 495 422 496
rect 422 495 423 496
rect 423 495 424 496
rect 424 495 425 496
rect 425 495 426 496
rect 426 495 427 496
rect 427 495 428 496
rect 428 495 429 496
rect 429 495 430 496
rect 430 495 431 496
rect 431 495 432 496
rect 432 495 433 496
rect 433 495 434 496
rect 434 495 435 496
rect 435 495 436 496
rect 436 495 437 496
rect 437 495 438 496
rect 438 495 439 496
rect 439 495 440 496
rect 440 495 441 496
rect 441 495 442 496
rect 442 495 443 496
rect 231 494 232 495
rect 232 494 233 495
rect 233 494 234 495
rect 234 494 235 495
rect 235 494 236 495
rect 236 494 237 495
rect 321 494 322 495
rect 322 494 323 495
rect 323 494 324 495
rect 324 494 325 495
rect 325 494 326 495
rect 326 494 327 495
rect 327 494 328 495
rect 328 494 329 495
rect 329 494 330 495
rect 330 494 331 495
rect 331 494 332 495
rect 332 494 333 495
rect 333 494 334 495
rect 334 494 335 495
rect 383 494 384 495
rect 384 494 385 495
rect 385 494 386 495
rect 386 494 387 495
rect 387 494 388 495
rect 388 494 389 495
rect 389 494 390 495
rect 390 494 391 495
rect 391 494 392 495
rect 392 494 393 495
rect 393 494 394 495
rect 394 494 395 495
rect 395 494 396 495
rect 396 494 397 495
rect 397 494 398 495
rect 412 494 413 495
rect 413 494 414 495
rect 414 494 415 495
rect 415 494 416 495
rect 416 494 417 495
rect 417 494 418 495
rect 418 494 419 495
rect 419 494 420 495
rect 420 494 421 495
rect 421 494 422 495
rect 422 494 423 495
rect 423 494 424 495
rect 424 494 425 495
rect 425 494 426 495
rect 426 494 427 495
rect 427 494 428 495
rect 428 494 429 495
rect 429 494 430 495
rect 430 494 431 495
rect 431 494 432 495
rect 432 494 433 495
rect 433 494 434 495
rect 434 494 435 495
rect 435 494 436 495
rect 436 494 437 495
rect 437 494 438 495
rect 438 494 439 495
rect 439 494 440 495
rect 440 494 441 495
rect 441 494 442 495
rect 442 494 443 495
rect 229 493 230 494
rect 230 493 231 494
rect 231 493 232 494
rect 232 493 233 494
rect 233 493 234 494
rect 234 493 235 494
rect 235 493 236 494
rect 236 493 237 494
rect 321 493 322 494
rect 322 493 323 494
rect 323 493 324 494
rect 324 493 325 494
rect 325 493 326 494
rect 326 493 327 494
rect 327 493 328 494
rect 328 493 329 494
rect 329 493 330 494
rect 330 493 331 494
rect 331 493 332 494
rect 332 493 333 494
rect 333 493 334 494
rect 334 493 335 494
rect 335 493 336 494
rect 336 493 337 494
rect 381 493 382 494
rect 382 493 383 494
rect 383 493 384 494
rect 384 493 385 494
rect 385 493 386 494
rect 386 493 387 494
rect 387 493 388 494
rect 388 493 389 494
rect 389 493 390 494
rect 390 493 391 494
rect 391 493 392 494
rect 392 493 393 494
rect 393 493 394 494
rect 394 493 395 494
rect 395 493 396 494
rect 396 493 397 494
rect 397 493 398 494
rect 412 493 413 494
rect 413 493 414 494
rect 414 493 415 494
rect 415 493 416 494
rect 416 493 417 494
rect 417 493 418 494
rect 418 493 419 494
rect 419 493 420 494
rect 420 493 421 494
rect 421 493 422 494
rect 422 493 423 494
rect 423 493 424 494
rect 424 493 425 494
rect 425 493 426 494
rect 426 493 427 494
rect 427 493 428 494
rect 428 493 429 494
rect 429 493 430 494
rect 430 493 431 494
rect 431 493 432 494
rect 432 493 433 494
rect 433 493 434 494
rect 434 493 435 494
rect 435 493 436 494
rect 436 493 437 494
rect 437 493 438 494
rect 438 493 439 494
rect 439 493 440 494
rect 440 493 441 494
rect 441 493 442 494
rect 442 493 443 494
rect 229 492 230 493
rect 230 492 231 493
rect 231 492 232 493
rect 232 492 233 493
rect 233 492 234 493
rect 324 492 325 493
rect 325 492 326 493
rect 326 492 327 493
rect 327 492 328 493
rect 328 492 329 493
rect 329 492 330 493
rect 330 492 331 493
rect 331 492 332 493
rect 332 492 333 493
rect 333 492 334 493
rect 334 492 335 493
rect 335 492 336 493
rect 336 492 337 493
rect 381 492 382 493
rect 382 492 383 493
rect 383 492 384 493
rect 384 492 385 493
rect 385 492 386 493
rect 386 492 387 493
rect 387 492 388 493
rect 388 492 389 493
rect 389 492 390 493
rect 390 492 391 493
rect 391 492 392 493
rect 392 492 393 493
rect 393 492 394 493
rect 394 492 395 493
rect 395 492 396 493
rect 396 492 397 493
rect 412 492 413 493
rect 413 492 414 493
rect 414 492 415 493
rect 415 492 416 493
rect 416 492 417 493
rect 417 492 418 493
rect 418 492 419 493
rect 419 492 420 493
rect 420 492 421 493
rect 421 492 422 493
rect 422 492 423 493
rect 423 492 424 493
rect 424 492 425 493
rect 425 492 426 493
rect 426 492 427 493
rect 427 492 428 493
rect 428 492 429 493
rect 429 492 430 493
rect 430 492 431 493
rect 431 492 432 493
rect 432 492 433 493
rect 433 492 434 493
rect 434 492 435 493
rect 435 492 436 493
rect 436 492 437 493
rect 437 492 438 493
rect 438 492 439 493
rect 439 492 440 493
rect 440 492 441 493
rect 441 492 442 493
rect 229 491 230 492
rect 230 491 231 492
rect 231 491 232 492
rect 232 491 233 492
rect 233 491 234 492
rect 324 491 325 492
rect 325 491 326 492
rect 326 491 327 492
rect 327 491 328 492
rect 328 491 329 492
rect 329 491 330 492
rect 330 491 331 492
rect 331 491 332 492
rect 332 491 333 492
rect 333 491 334 492
rect 334 491 335 492
rect 335 491 336 492
rect 336 491 337 492
rect 337 491 338 492
rect 338 491 339 492
rect 379 491 380 492
rect 380 491 381 492
rect 381 491 382 492
rect 382 491 383 492
rect 383 491 384 492
rect 384 491 385 492
rect 385 491 386 492
rect 386 491 387 492
rect 387 491 388 492
rect 388 491 389 492
rect 389 491 390 492
rect 390 491 391 492
rect 391 491 392 492
rect 392 491 393 492
rect 393 491 394 492
rect 394 491 395 492
rect 395 491 396 492
rect 396 491 397 492
rect 412 491 413 492
rect 413 491 414 492
rect 414 491 415 492
rect 415 491 416 492
rect 416 491 417 492
rect 417 491 418 492
rect 418 491 419 492
rect 419 491 420 492
rect 420 491 421 492
rect 421 491 422 492
rect 422 491 423 492
rect 423 491 424 492
rect 424 491 425 492
rect 425 491 426 492
rect 426 491 427 492
rect 427 491 428 492
rect 428 491 429 492
rect 429 491 430 492
rect 430 491 431 492
rect 431 491 432 492
rect 432 491 433 492
rect 433 491 434 492
rect 434 491 435 492
rect 435 491 436 492
rect 436 491 437 492
rect 437 491 438 492
rect 438 491 439 492
rect 439 491 440 492
rect 440 491 441 492
rect 441 491 442 492
rect 442 491 443 492
rect 328 490 329 491
rect 329 490 330 491
rect 330 490 331 491
rect 331 490 332 491
rect 332 490 333 491
rect 333 490 334 491
rect 334 490 335 491
rect 335 490 336 491
rect 336 490 337 491
rect 337 490 338 491
rect 338 490 339 491
rect 379 490 380 491
rect 380 490 381 491
rect 381 490 382 491
rect 382 490 383 491
rect 383 490 384 491
rect 384 490 385 491
rect 385 490 386 491
rect 386 490 387 491
rect 387 490 388 491
rect 388 490 389 491
rect 389 490 390 491
rect 390 490 391 491
rect 391 490 392 491
rect 392 490 393 491
rect 412 490 413 491
rect 413 490 414 491
rect 414 490 415 491
rect 415 490 416 491
rect 416 490 417 491
rect 417 490 418 491
rect 418 490 419 491
rect 419 490 420 491
rect 420 490 421 491
rect 421 490 422 491
rect 422 490 423 491
rect 423 490 424 491
rect 424 490 425 491
rect 425 490 426 491
rect 426 490 427 491
rect 427 490 428 491
rect 428 490 429 491
rect 429 490 430 491
rect 430 490 431 491
rect 431 490 432 491
rect 432 490 433 491
rect 433 490 434 491
rect 434 490 435 491
rect 435 490 436 491
rect 436 490 437 491
rect 437 490 438 491
rect 438 490 439 491
rect 439 490 440 491
rect 440 490 441 491
rect 441 490 442 491
rect 442 490 443 491
rect 328 489 329 490
rect 329 489 330 490
rect 330 489 331 490
rect 331 489 332 490
rect 332 489 333 490
rect 333 489 334 490
rect 334 489 335 490
rect 335 489 336 490
rect 336 489 337 490
rect 337 489 338 490
rect 338 489 339 490
rect 339 489 340 490
rect 340 489 341 490
rect 341 489 342 490
rect 377 489 378 490
rect 378 489 379 490
rect 379 489 380 490
rect 380 489 381 490
rect 381 489 382 490
rect 382 489 383 490
rect 383 489 384 490
rect 384 489 385 490
rect 385 489 386 490
rect 386 489 387 490
rect 387 489 388 490
rect 388 489 389 490
rect 389 489 390 490
rect 390 489 391 490
rect 391 489 392 490
rect 392 489 393 490
rect 412 489 413 490
rect 413 489 414 490
rect 414 489 415 490
rect 415 489 416 490
rect 416 489 417 490
rect 417 489 418 490
rect 418 489 419 490
rect 419 489 420 490
rect 420 489 421 490
rect 421 489 422 490
rect 422 489 423 490
rect 423 489 424 490
rect 424 489 425 490
rect 425 489 426 490
rect 426 489 427 490
rect 427 489 428 490
rect 428 489 429 490
rect 429 489 430 490
rect 430 489 431 490
rect 431 489 432 490
rect 432 489 433 490
rect 433 489 434 490
rect 434 489 435 490
rect 435 489 436 490
rect 436 489 437 490
rect 437 489 438 490
rect 438 489 439 490
rect 439 489 440 490
rect 440 489 441 490
rect 441 489 442 490
rect 442 489 443 490
rect 330 488 331 489
rect 331 488 332 489
rect 332 488 333 489
rect 333 488 334 489
rect 334 488 335 489
rect 335 488 336 489
rect 336 488 337 489
rect 337 488 338 489
rect 338 488 339 489
rect 339 488 340 489
rect 340 488 341 489
rect 341 488 342 489
rect 377 488 378 489
rect 378 488 379 489
rect 379 488 380 489
rect 380 488 381 489
rect 381 488 382 489
rect 382 488 383 489
rect 383 488 384 489
rect 384 488 385 489
rect 385 488 386 489
rect 386 488 387 489
rect 387 488 388 489
rect 388 488 389 489
rect 389 488 390 489
rect 390 488 391 489
rect 412 488 413 489
rect 413 488 414 489
rect 414 488 415 489
rect 415 488 416 489
rect 416 488 417 489
rect 417 488 418 489
rect 418 488 419 489
rect 419 488 420 489
rect 420 488 421 489
rect 421 488 422 489
rect 422 488 423 489
rect 423 488 424 489
rect 424 488 425 489
rect 425 488 426 489
rect 426 488 427 489
rect 427 488 428 489
rect 428 488 429 489
rect 429 488 430 489
rect 430 488 431 489
rect 431 488 432 489
rect 432 488 433 489
rect 433 488 434 489
rect 434 488 435 489
rect 435 488 436 489
rect 436 488 437 489
rect 437 488 438 489
rect 438 488 439 489
rect 439 488 440 489
rect 440 488 441 489
rect 441 488 442 489
rect 442 488 443 489
rect 221 487 222 488
rect 222 487 223 488
rect 223 487 224 488
rect 330 487 331 488
rect 331 487 332 488
rect 332 487 333 488
rect 333 487 334 488
rect 334 487 335 488
rect 335 487 336 488
rect 336 487 337 488
rect 337 487 338 488
rect 338 487 339 488
rect 339 487 340 488
rect 340 487 341 488
rect 341 487 342 488
rect 342 487 343 488
rect 343 487 344 488
rect 375 487 376 488
rect 376 487 377 488
rect 377 487 378 488
rect 378 487 379 488
rect 379 487 380 488
rect 380 487 381 488
rect 381 487 382 488
rect 382 487 383 488
rect 383 487 384 488
rect 384 487 385 488
rect 385 487 386 488
rect 386 487 387 488
rect 387 487 388 488
rect 388 487 389 488
rect 389 487 390 488
rect 390 487 391 488
rect 412 487 413 488
rect 413 487 414 488
rect 414 487 415 488
rect 415 487 416 488
rect 416 487 417 488
rect 417 487 418 488
rect 418 487 419 488
rect 419 487 420 488
rect 420 487 421 488
rect 421 487 422 488
rect 422 487 423 488
rect 423 487 424 488
rect 424 487 425 488
rect 425 487 426 488
rect 426 487 427 488
rect 427 487 428 488
rect 428 487 429 488
rect 429 487 430 488
rect 430 487 431 488
rect 431 487 432 488
rect 432 487 433 488
rect 433 487 434 488
rect 434 487 435 488
rect 435 487 436 488
rect 436 487 437 488
rect 437 487 438 488
rect 438 487 439 488
rect 439 487 440 488
rect 440 487 441 488
rect 441 487 442 488
rect 442 487 443 488
rect 221 486 222 487
rect 222 486 223 487
rect 223 486 224 487
rect 334 486 335 487
rect 335 486 336 487
rect 336 486 337 487
rect 337 486 338 487
rect 338 486 339 487
rect 339 486 340 487
rect 340 486 341 487
rect 341 486 342 487
rect 342 486 343 487
rect 343 486 344 487
rect 375 486 376 487
rect 376 486 377 487
rect 377 486 378 487
rect 378 486 379 487
rect 379 486 380 487
rect 380 486 381 487
rect 381 486 382 487
rect 382 486 383 487
rect 383 486 384 487
rect 384 486 385 487
rect 385 486 386 487
rect 386 486 387 487
rect 387 486 388 487
rect 388 486 389 487
rect 414 486 415 487
rect 415 486 416 487
rect 416 486 417 487
rect 417 486 418 487
rect 418 486 419 487
rect 419 486 420 487
rect 420 486 421 487
rect 421 486 422 487
rect 422 486 423 487
rect 423 486 424 487
rect 424 486 425 487
rect 425 486 426 487
rect 426 486 427 487
rect 427 486 428 487
rect 428 486 429 487
rect 429 486 430 487
rect 430 486 431 487
rect 431 486 432 487
rect 432 486 433 487
rect 433 486 434 487
rect 434 486 435 487
rect 435 486 436 487
rect 436 486 437 487
rect 437 486 438 487
rect 438 486 439 487
rect 439 486 440 487
rect 440 486 441 487
rect 441 486 442 487
rect 220 485 221 486
rect 221 485 222 486
rect 222 485 223 486
rect 223 485 224 486
rect 334 485 335 486
rect 335 485 336 486
rect 336 485 337 486
rect 337 485 338 486
rect 338 485 339 486
rect 339 485 340 486
rect 340 485 341 486
rect 341 485 342 486
rect 342 485 343 486
rect 343 485 344 486
rect 344 485 345 486
rect 345 485 346 486
rect 373 485 374 486
rect 374 485 375 486
rect 375 485 376 486
rect 376 485 377 486
rect 377 485 378 486
rect 378 485 379 486
rect 379 485 380 486
rect 380 485 381 486
rect 381 485 382 486
rect 382 485 383 486
rect 383 485 384 486
rect 384 485 385 486
rect 385 485 386 486
rect 386 485 387 486
rect 387 485 388 486
rect 388 485 389 486
rect 412 485 413 486
rect 413 485 414 486
rect 414 485 415 486
rect 415 485 416 486
rect 416 485 417 486
rect 417 485 418 486
rect 418 485 419 486
rect 419 485 420 486
rect 420 485 421 486
rect 421 485 422 486
rect 422 485 423 486
rect 423 485 424 486
rect 424 485 425 486
rect 425 485 426 486
rect 426 485 427 486
rect 427 485 428 486
rect 428 485 429 486
rect 429 485 430 486
rect 430 485 431 486
rect 431 485 432 486
rect 432 485 433 486
rect 433 485 434 486
rect 434 485 435 486
rect 435 485 436 486
rect 436 485 437 486
rect 437 485 438 486
rect 438 485 439 486
rect 439 485 440 486
rect 440 485 441 486
rect 441 485 442 486
rect 442 485 443 486
rect 220 484 221 485
rect 221 484 222 485
rect 336 484 337 485
rect 337 484 338 485
rect 338 484 339 485
rect 339 484 340 485
rect 340 484 341 485
rect 341 484 342 485
rect 342 484 343 485
rect 343 484 344 485
rect 344 484 345 485
rect 345 484 346 485
rect 373 484 374 485
rect 374 484 375 485
rect 375 484 376 485
rect 376 484 377 485
rect 377 484 378 485
rect 378 484 379 485
rect 379 484 380 485
rect 380 484 381 485
rect 381 484 382 485
rect 382 484 383 485
rect 383 484 384 485
rect 384 484 385 485
rect 385 484 386 485
rect 386 484 387 485
rect 412 484 413 485
rect 413 484 414 485
rect 414 484 415 485
rect 415 484 416 485
rect 416 484 417 485
rect 417 484 418 485
rect 418 484 419 485
rect 419 484 420 485
rect 420 484 421 485
rect 421 484 422 485
rect 422 484 423 485
rect 423 484 424 485
rect 424 484 425 485
rect 425 484 426 485
rect 426 484 427 485
rect 427 484 428 485
rect 428 484 429 485
rect 429 484 430 485
rect 430 484 431 485
rect 431 484 432 485
rect 432 484 433 485
rect 433 484 434 485
rect 434 484 435 485
rect 435 484 436 485
rect 436 484 437 485
rect 437 484 438 485
rect 438 484 439 485
rect 439 484 440 485
rect 440 484 441 485
rect 441 484 442 485
rect 442 484 443 485
rect 220 483 221 484
rect 221 483 222 484
rect 336 483 337 484
rect 337 483 338 484
rect 338 483 339 484
rect 339 483 340 484
rect 340 483 341 484
rect 341 483 342 484
rect 342 483 343 484
rect 343 483 344 484
rect 344 483 345 484
rect 345 483 346 484
rect 373 483 374 484
rect 374 483 375 484
rect 375 483 376 484
rect 376 483 377 484
rect 377 483 378 484
rect 378 483 379 484
rect 379 483 380 484
rect 380 483 381 484
rect 381 483 382 484
rect 382 483 383 484
rect 383 483 384 484
rect 384 483 385 484
rect 385 483 386 484
rect 386 483 387 484
rect 412 483 413 484
rect 413 483 414 484
rect 414 483 415 484
rect 415 483 416 484
rect 416 483 417 484
rect 417 483 418 484
rect 418 483 419 484
rect 419 483 420 484
rect 420 483 421 484
rect 421 483 422 484
rect 422 483 423 484
rect 423 483 424 484
rect 424 483 425 484
rect 425 483 426 484
rect 426 483 427 484
rect 427 483 428 484
rect 428 483 429 484
rect 429 483 430 484
rect 430 483 431 484
rect 431 483 432 484
rect 432 483 433 484
rect 433 483 434 484
rect 434 483 435 484
rect 435 483 436 484
rect 436 483 437 484
rect 437 483 438 484
rect 438 483 439 484
rect 439 483 440 484
rect 440 483 441 484
rect 441 483 442 484
rect 442 483 443 484
rect 218 482 219 483
rect 219 482 220 483
rect 220 482 221 483
rect 221 482 222 483
rect 336 482 337 483
rect 337 482 338 483
rect 338 482 339 483
rect 339 482 340 483
rect 340 482 341 483
rect 341 482 342 483
rect 342 482 343 483
rect 343 482 344 483
rect 344 482 345 483
rect 345 482 346 483
rect 346 482 347 483
rect 347 482 348 483
rect 371 482 372 483
rect 372 482 373 483
rect 373 482 374 483
rect 374 482 375 483
rect 375 482 376 483
rect 376 482 377 483
rect 377 482 378 483
rect 378 482 379 483
rect 379 482 380 483
rect 380 482 381 483
rect 381 482 382 483
rect 382 482 383 483
rect 383 482 384 483
rect 384 482 385 483
rect 385 482 386 483
rect 386 482 387 483
rect 412 482 413 483
rect 413 482 414 483
rect 414 482 415 483
rect 415 482 416 483
rect 416 482 417 483
rect 417 482 418 483
rect 418 482 419 483
rect 419 482 420 483
rect 420 482 421 483
rect 421 482 422 483
rect 422 482 423 483
rect 423 482 424 483
rect 424 482 425 483
rect 425 482 426 483
rect 426 482 427 483
rect 427 482 428 483
rect 428 482 429 483
rect 429 482 430 483
rect 430 482 431 483
rect 431 482 432 483
rect 432 482 433 483
rect 433 482 434 483
rect 434 482 435 483
rect 435 482 436 483
rect 436 482 437 483
rect 437 482 438 483
rect 438 482 439 483
rect 439 482 440 483
rect 440 482 441 483
rect 441 482 442 483
rect 442 482 443 483
rect 218 481 219 482
rect 219 481 220 482
rect 220 481 221 482
rect 338 481 339 482
rect 339 481 340 482
rect 340 481 341 482
rect 341 481 342 482
rect 342 481 343 482
rect 343 481 344 482
rect 344 481 345 482
rect 345 481 346 482
rect 346 481 347 482
rect 347 481 348 482
rect 371 481 372 482
rect 372 481 373 482
rect 373 481 374 482
rect 374 481 375 482
rect 375 481 376 482
rect 376 481 377 482
rect 377 481 378 482
rect 378 481 379 482
rect 379 481 380 482
rect 380 481 381 482
rect 381 481 382 482
rect 382 481 383 482
rect 383 481 384 482
rect 384 481 385 482
rect 412 481 413 482
rect 413 481 414 482
rect 414 481 415 482
rect 415 481 416 482
rect 416 481 417 482
rect 417 481 418 482
rect 418 481 419 482
rect 419 481 420 482
rect 420 481 421 482
rect 421 481 422 482
rect 422 481 423 482
rect 423 481 424 482
rect 424 481 425 482
rect 425 481 426 482
rect 426 481 427 482
rect 427 481 428 482
rect 428 481 429 482
rect 429 481 430 482
rect 430 481 431 482
rect 431 481 432 482
rect 432 481 433 482
rect 433 481 434 482
rect 434 481 435 482
rect 435 481 436 482
rect 436 481 437 482
rect 437 481 438 482
rect 438 481 439 482
rect 439 481 440 482
rect 440 481 441 482
rect 441 481 442 482
rect 442 481 443 482
rect 214 480 215 481
rect 215 480 216 481
rect 216 480 217 481
rect 217 480 218 481
rect 218 480 219 481
rect 219 480 220 481
rect 220 480 221 481
rect 338 480 339 481
rect 339 480 340 481
rect 340 480 341 481
rect 341 480 342 481
rect 342 480 343 481
rect 343 480 344 481
rect 344 480 345 481
rect 345 480 346 481
rect 346 480 347 481
rect 347 480 348 481
rect 348 480 349 481
rect 349 480 350 481
rect 350 480 351 481
rect 351 480 352 481
rect 369 480 370 481
rect 370 480 371 481
rect 371 480 372 481
rect 372 480 373 481
rect 373 480 374 481
rect 374 480 375 481
rect 375 480 376 481
rect 376 480 377 481
rect 377 480 378 481
rect 378 480 379 481
rect 379 480 380 481
rect 380 480 381 481
rect 381 480 382 481
rect 382 480 383 481
rect 383 480 384 481
rect 384 480 385 481
rect 412 480 413 481
rect 413 480 414 481
rect 414 480 415 481
rect 415 480 416 481
rect 416 480 417 481
rect 417 480 418 481
rect 418 480 419 481
rect 419 480 420 481
rect 420 480 421 481
rect 421 480 422 481
rect 422 480 423 481
rect 423 480 424 481
rect 424 480 425 481
rect 425 480 426 481
rect 426 480 427 481
rect 427 480 428 481
rect 428 480 429 481
rect 429 480 430 481
rect 430 480 431 481
rect 431 480 432 481
rect 432 480 433 481
rect 433 480 434 481
rect 434 480 435 481
rect 435 480 436 481
rect 436 480 437 481
rect 437 480 438 481
rect 438 480 439 481
rect 439 480 440 481
rect 440 480 441 481
rect 441 480 442 481
rect 442 480 443 481
rect 214 479 215 480
rect 215 479 216 480
rect 216 479 217 480
rect 217 479 218 480
rect 218 479 219 480
rect 339 479 340 480
rect 340 479 341 480
rect 341 479 342 480
rect 342 479 343 480
rect 343 479 344 480
rect 344 479 345 480
rect 345 479 346 480
rect 346 479 347 480
rect 347 479 348 480
rect 348 479 349 480
rect 349 479 350 480
rect 350 479 351 480
rect 351 479 352 480
rect 369 479 370 480
rect 370 479 371 480
rect 371 479 372 480
rect 372 479 373 480
rect 373 479 374 480
rect 374 479 375 480
rect 375 479 376 480
rect 376 479 377 480
rect 377 479 378 480
rect 378 479 379 480
rect 379 479 380 480
rect 380 479 381 480
rect 381 479 382 480
rect 382 479 383 480
rect 383 479 384 480
rect 412 479 413 480
rect 413 479 414 480
rect 414 479 415 480
rect 415 479 416 480
rect 416 479 417 480
rect 417 479 418 480
rect 418 479 419 480
rect 419 479 420 480
rect 420 479 421 480
rect 421 479 422 480
rect 422 479 423 480
rect 423 479 424 480
rect 424 479 425 480
rect 425 479 426 480
rect 426 479 427 480
rect 427 479 428 480
rect 428 479 429 480
rect 429 479 430 480
rect 430 479 431 480
rect 431 479 432 480
rect 432 479 433 480
rect 433 479 434 480
rect 434 479 435 480
rect 435 479 436 480
rect 436 479 437 480
rect 437 479 438 480
rect 438 479 439 480
rect 439 479 440 480
rect 440 479 441 480
rect 441 479 442 480
rect 442 479 443 480
rect 214 478 215 479
rect 215 478 216 479
rect 216 478 217 479
rect 217 478 218 479
rect 218 478 219 479
rect 339 478 340 479
rect 340 478 341 479
rect 341 478 342 479
rect 342 478 343 479
rect 343 478 344 479
rect 344 478 345 479
rect 345 478 346 479
rect 346 478 347 479
rect 347 478 348 479
rect 348 478 349 479
rect 349 478 350 479
rect 350 478 351 479
rect 351 478 352 479
rect 352 478 353 479
rect 353 478 354 479
rect 366 478 367 479
rect 367 478 368 479
rect 368 478 369 479
rect 369 478 370 479
rect 370 478 371 479
rect 371 478 372 479
rect 372 478 373 479
rect 373 478 374 479
rect 374 478 375 479
rect 375 478 376 479
rect 376 478 377 479
rect 377 478 378 479
rect 378 478 379 479
rect 379 478 380 479
rect 380 478 381 479
rect 381 478 382 479
rect 382 478 383 479
rect 383 478 384 479
rect 412 478 413 479
rect 413 478 414 479
rect 414 478 415 479
rect 415 478 416 479
rect 416 478 417 479
rect 417 478 418 479
rect 418 478 419 479
rect 419 478 420 479
rect 420 478 421 479
rect 421 478 422 479
rect 422 478 423 479
rect 423 478 424 479
rect 424 478 425 479
rect 425 478 426 479
rect 426 478 427 479
rect 427 478 428 479
rect 428 478 429 479
rect 429 478 430 479
rect 430 478 431 479
rect 431 478 432 479
rect 432 478 433 479
rect 433 478 434 479
rect 434 478 435 479
rect 435 478 436 479
rect 436 478 437 479
rect 437 478 438 479
rect 438 478 439 479
rect 439 478 440 479
rect 440 478 441 479
rect 441 478 442 479
rect 442 478 443 479
rect 214 477 215 478
rect 215 477 216 478
rect 216 477 217 478
rect 341 477 342 478
rect 342 477 343 478
rect 343 477 344 478
rect 344 477 345 478
rect 345 477 346 478
rect 346 477 347 478
rect 347 477 348 478
rect 348 477 349 478
rect 349 477 350 478
rect 350 477 351 478
rect 351 477 352 478
rect 352 477 353 478
rect 353 477 354 478
rect 366 477 367 478
rect 367 477 368 478
rect 368 477 369 478
rect 369 477 370 478
rect 370 477 371 478
rect 371 477 372 478
rect 372 477 373 478
rect 373 477 374 478
rect 374 477 375 478
rect 375 477 376 478
rect 376 477 377 478
rect 377 477 378 478
rect 378 477 379 478
rect 379 477 380 478
rect 380 477 381 478
rect 381 477 382 478
rect 412 477 413 478
rect 413 477 414 478
rect 414 477 415 478
rect 415 477 416 478
rect 416 477 417 478
rect 417 477 418 478
rect 418 477 419 478
rect 419 477 420 478
rect 420 477 421 478
rect 421 477 422 478
rect 422 477 423 478
rect 423 477 424 478
rect 424 477 425 478
rect 425 477 426 478
rect 426 477 427 478
rect 427 477 428 478
rect 428 477 429 478
rect 429 477 430 478
rect 430 477 431 478
rect 431 477 432 478
rect 432 477 433 478
rect 433 477 434 478
rect 434 477 435 478
rect 435 477 436 478
rect 436 477 437 478
rect 437 477 438 478
rect 438 477 439 478
rect 439 477 440 478
rect 212 476 213 477
rect 213 476 214 477
rect 214 476 215 477
rect 215 476 216 477
rect 216 476 217 477
rect 341 476 342 477
rect 342 476 343 477
rect 343 476 344 477
rect 344 476 345 477
rect 345 476 346 477
rect 346 476 347 477
rect 347 476 348 477
rect 348 476 349 477
rect 349 476 350 477
rect 350 476 351 477
rect 351 476 352 477
rect 352 476 353 477
rect 353 476 354 477
rect 354 476 355 477
rect 364 476 365 477
rect 365 476 366 477
rect 366 476 367 477
rect 367 476 368 477
rect 368 476 369 477
rect 369 476 370 477
rect 370 476 371 477
rect 371 476 372 477
rect 372 476 373 477
rect 373 476 374 477
rect 374 476 375 477
rect 375 476 376 477
rect 376 476 377 477
rect 377 476 378 477
rect 378 476 379 477
rect 379 476 380 477
rect 380 476 381 477
rect 381 476 382 477
rect 412 476 413 477
rect 413 476 414 477
rect 414 476 415 477
rect 415 476 416 477
rect 416 476 417 477
rect 417 476 418 477
rect 418 476 419 477
rect 419 476 420 477
rect 420 476 421 477
rect 421 476 422 477
rect 422 476 423 477
rect 423 476 424 477
rect 424 476 425 477
rect 425 476 426 477
rect 426 476 427 477
rect 427 476 428 477
rect 428 476 429 477
rect 429 476 430 477
rect 430 476 431 477
rect 431 476 432 477
rect 432 476 433 477
rect 433 476 434 477
rect 434 476 435 477
rect 435 476 436 477
rect 436 476 437 477
rect 437 476 438 477
rect 438 476 439 477
rect 439 476 440 477
rect 212 475 213 476
rect 213 475 214 476
rect 214 475 215 476
rect 343 475 344 476
rect 344 475 345 476
rect 345 475 346 476
rect 346 475 347 476
rect 347 475 348 476
rect 348 475 349 476
rect 349 475 350 476
rect 350 475 351 476
rect 351 475 352 476
rect 352 475 353 476
rect 353 475 354 476
rect 354 475 355 476
rect 364 475 365 476
rect 365 475 366 476
rect 366 475 367 476
rect 367 475 368 476
rect 368 475 369 476
rect 369 475 370 476
rect 370 475 371 476
rect 371 475 372 476
rect 372 475 373 476
rect 373 475 374 476
rect 374 475 375 476
rect 375 475 376 476
rect 376 475 377 476
rect 377 475 378 476
rect 378 475 379 476
rect 379 475 380 476
rect 412 475 413 476
rect 413 475 414 476
rect 414 475 415 476
rect 415 475 416 476
rect 416 475 417 476
rect 417 475 418 476
rect 418 475 419 476
rect 419 475 420 476
rect 420 475 421 476
rect 421 475 422 476
rect 422 475 423 476
rect 423 475 424 476
rect 424 475 425 476
rect 425 475 426 476
rect 426 475 427 476
rect 427 475 428 476
rect 428 475 429 476
rect 429 475 430 476
rect 430 475 431 476
rect 431 475 432 476
rect 432 475 433 476
rect 433 475 434 476
rect 434 475 435 476
rect 435 475 436 476
rect 210 474 211 475
rect 211 474 212 475
rect 212 474 213 475
rect 213 474 214 475
rect 214 474 215 475
rect 343 474 344 475
rect 344 474 345 475
rect 345 474 346 475
rect 346 474 347 475
rect 347 474 348 475
rect 348 474 349 475
rect 349 474 350 475
rect 350 474 351 475
rect 351 474 352 475
rect 352 474 353 475
rect 353 474 354 475
rect 354 474 355 475
rect 355 474 356 475
rect 356 474 357 475
rect 357 474 358 475
rect 358 474 359 475
rect 360 474 361 475
rect 361 474 362 475
rect 362 474 363 475
rect 363 474 364 475
rect 364 474 365 475
rect 365 474 366 475
rect 366 474 367 475
rect 367 474 368 475
rect 368 474 369 475
rect 369 474 370 475
rect 370 474 371 475
rect 371 474 372 475
rect 372 474 373 475
rect 373 474 374 475
rect 374 474 375 475
rect 375 474 376 475
rect 376 474 377 475
rect 377 474 378 475
rect 378 474 379 475
rect 379 474 380 475
rect 412 474 413 475
rect 413 474 414 475
rect 414 474 415 475
rect 415 474 416 475
rect 416 474 417 475
rect 417 474 418 475
rect 418 474 419 475
rect 419 474 420 475
rect 420 474 421 475
rect 421 474 422 475
rect 422 474 423 475
rect 423 474 424 475
rect 424 474 425 475
rect 425 474 426 475
rect 426 474 427 475
rect 427 474 428 475
rect 428 474 429 475
rect 429 474 430 475
rect 430 474 431 475
rect 431 474 432 475
rect 432 474 433 475
rect 433 474 434 475
rect 434 474 435 475
rect 435 474 436 475
rect 210 473 211 474
rect 211 473 212 474
rect 212 473 213 474
rect 213 473 214 474
rect 214 473 215 474
rect 345 473 346 474
rect 346 473 347 474
rect 347 473 348 474
rect 348 473 349 474
rect 349 473 350 474
rect 350 473 351 474
rect 351 473 352 474
rect 352 473 353 474
rect 353 473 354 474
rect 354 473 355 474
rect 355 473 356 474
rect 356 473 357 474
rect 357 473 358 474
rect 358 473 359 474
rect 360 473 361 474
rect 361 473 362 474
rect 362 473 363 474
rect 363 473 364 474
rect 364 473 365 474
rect 365 473 366 474
rect 366 473 367 474
rect 367 473 368 474
rect 368 473 369 474
rect 369 473 370 474
rect 370 473 371 474
rect 371 473 372 474
rect 372 473 373 474
rect 373 473 374 474
rect 374 473 375 474
rect 375 473 376 474
rect 376 473 377 474
rect 377 473 378 474
rect 378 473 379 474
rect 379 473 380 474
rect 412 473 413 474
rect 413 473 414 474
rect 414 473 415 474
rect 415 473 416 474
rect 416 473 417 474
rect 417 473 418 474
rect 418 473 419 474
rect 419 473 420 474
rect 420 473 421 474
rect 421 473 422 474
rect 422 473 423 474
rect 423 473 424 474
rect 424 473 425 474
rect 425 473 426 474
rect 426 473 427 474
rect 427 473 428 474
rect 428 473 429 474
rect 429 473 430 474
rect 208 472 209 473
rect 209 472 210 473
rect 210 472 211 473
rect 211 472 212 473
rect 212 472 213 473
rect 213 472 214 473
rect 214 472 215 473
rect 345 472 346 473
rect 346 472 347 473
rect 347 472 348 473
rect 348 472 349 473
rect 349 472 350 473
rect 350 472 351 473
rect 351 472 352 473
rect 352 472 353 473
rect 353 472 354 473
rect 354 472 355 473
rect 355 472 356 473
rect 356 472 357 473
rect 357 472 358 473
rect 358 472 359 473
rect 359 472 360 473
rect 360 472 361 473
rect 361 472 362 473
rect 362 472 363 473
rect 363 472 364 473
rect 364 472 365 473
rect 365 472 366 473
rect 366 472 367 473
rect 367 472 368 473
rect 368 472 369 473
rect 369 472 370 473
rect 370 472 371 473
rect 371 472 372 473
rect 372 472 373 473
rect 373 472 374 473
rect 374 472 375 473
rect 375 472 376 473
rect 376 472 377 473
rect 377 472 378 473
rect 378 472 379 473
rect 379 472 380 473
rect 411 472 412 473
rect 412 472 413 473
rect 413 472 414 473
rect 414 472 415 473
rect 415 472 416 473
rect 416 472 417 473
rect 417 472 418 473
rect 418 472 419 473
rect 419 472 420 473
rect 420 472 421 473
rect 421 472 422 473
rect 422 472 423 473
rect 423 472 424 473
rect 424 472 425 473
rect 425 472 426 473
rect 426 472 427 473
rect 427 472 428 473
rect 428 472 429 473
rect 429 472 430 473
rect 208 471 209 472
rect 209 471 210 472
rect 210 471 211 472
rect 345 471 346 472
rect 346 471 347 472
rect 347 471 348 472
rect 348 471 349 472
rect 349 471 350 472
rect 350 471 351 472
rect 351 471 352 472
rect 352 471 353 472
rect 353 471 354 472
rect 354 471 355 472
rect 355 471 356 472
rect 356 471 357 472
rect 357 471 358 472
rect 358 471 359 472
rect 359 471 360 472
rect 360 471 361 472
rect 361 471 362 472
rect 362 471 363 472
rect 363 471 364 472
rect 364 471 365 472
rect 365 471 366 472
rect 366 471 367 472
rect 367 471 368 472
rect 368 471 369 472
rect 369 471 370 472
rect 370 471 371 472
rect 371 471 372 472
rect 372 471 373 472
rect 373 471 374 472
rect 374 471 375 472
rect 375 471 376 472
rect 376 471 377 472
rect 377 471 378 472
rect 411 471 412 472
rect 412 471 413 472
rect 413 471 414 472
rect 414 471 415 472
rect 415 471 416 472
rect 416 471 417 472
rect 417 471 418 472
rect 418 471 419 472
rect 419 471 420 472
rect 420 471 421 472
rect 421 471 422 472
rect 422 471 423 472
rect 423 471 424 472
rect 424 471 425 472
rect 425 471 426 472
rect 426 471 427 472
rect 206 470 207 471
rect 207 470 208 471
rect 208 470 209 471
rect 209 470 210 471
rect 210 470 211 471
rect 345 470 346 471
rect 346 470 347 471
rect 347 470 348 471
rect 348 470 349 471
rect 349 470 350 471
rect 350 470 351 471
rect 351 470 352 471
rect 352 470 353 471
rect 353 470 354 471
rect 354 470 355 471
rect 355 470 356 471
rect 356 470 357 471
rect 357 470 358 471
rect 358 470 359 471
rect 359 470 360 471
rect 360 470 361 471
rect 361 470 362 471
rect 362 470 363 471
rect 363 470 364 471
rect 364 470 365 471
rect 365 470 366 471
rect 366 470 367 471
rect 367 470 368 471
rect 368 470 369 471
rect 369 470 370 471
rect 370 470 371 471
rect 371 470 372 471
rect 372 470 373 471
rect 373 470 374 471
rect 374 470 375 471
rect 375 470 376 471
rect 376 470 377 471
rect 377 470 378 471
rect 409 470 410 471
rect 410 470 411 471
rect 411 470 412 471
rect 412 470 413 471
rect 413 470 414 471
rect 414 470 415 471
rect 415 470 416 471
rect 416 470 417 471
rect 417 470 418 471
rect 418 470 419 471
rect 419 470 420 471
rect 420 470 421 471
rect 421 470 422 471
rect 422 470 423 471
rect 423 470 424 471
rect 424 470 425 471
rect 425 470 426 471
rect 426 470 427 471
rect 206 469 207 470
rect 207 469 208 470
rect 208 469 209 470
rect 347 469 348 470
rect 348 469 349 470
rect 349 469 350 470
rect 350 469 351 470
rect 351 469 352 470
rect 352 469 353 470
rect 353 469 354 470
rect 354 469 355 470
rect 355 469 356 470
rect 356 469 357 470
rect 357 469 358 470
rect 358 469 359 470
rect 359 469 360 470
rect 360 469 361 470
rect 361 469 362 470
rect 362 469 363 470
rect 363 469 364 470
rect 364 469 365 470
rect 365 469 366 470
rect 366 469 367 470
rect 367 469 368 470
rect 368 469 369 470
rect 369 469 370 470
rect 370 469 371 470
rect 371 469 372 470
rect 372 469 373 470
rect 373 469 374 470
rect 374 469 375 470
rect 375 469 376 470
rect 409 469 410 470
rect 410 469 411 470
rect 411 469 412 470
rect 412 469 413 470
rect 413 469 414 470
rect 414 469 415 470
rect 415 469 416 470
rect 416 469 417 470
rect 417 469 418 470
rect 418 469 419 470
rect 419 469 420 470
rect 420 469 421 470
rect 421 469 422 470
rect 422 469 423 470
rect 423 469 424 470
rect 424 469 425 470
rect 203 468 204 469
rect 204 468 205 469
rect 205 468 206 469
rect 206 468 207 469
rect 207 468 208 469
rect 208 468 209 469
rect 347 468 348 469
rect 348 468 349 469
rect 349 468 350 469
rect 350 468 351 469
rect 351 468 352 469
rect 352 468 353 469
rect 353 468 354 469
rect 354 468 355 469
rect 355 468 356 469
rect 356 468 357 469
rect 357 468 358 469
rect 358 468 359 469
rect 359 468 360 469
rect 360 468 361 469
rect 361 468 362 469
rect 362 468 363 469
rect 363 468 364 469
rect 364 468 365 469
rect 365 468 366 469
rect 366 468 367 469
rect 367 468 368 469
rect 368 468 369 469
rect 369 468 370 469
rect 370 468 371 469
rect 371 468 372 469
rect 372 468 373 469
rect 373 468 374 469
rect 374 468 375 469
rect 375 468 376 469
rect 409 468 410 469
rect 410 468 411 469
rect 411 468 412 469
rect 412 468 413 469
rect 413 468 414 469
rect 414 468 415 469
rect 415 468 416 469
rect 416 468 417 469
rect 417 468 418 469
rect 418 468 419 469
rect 419 468 420 469
rect 420 468 421 469
rect 421 468 422 469
rect 422 468 423 469
rect 423 468 424 469
rect 424 468 425 469
rect 203 467 204 468
rect 204 467 205 468
rect 205 467 206 468
rect 206 467 207 468
rect 207 467 208 468
rect 208 467 209 468
rect 347 467 348 468
rect 348 467 349 468
rect 349 467 350 468
rect 350 467 351 468
rect 351 467 352 468
rect 352 467 353 468
rect 353 467 354 468
rect 354 467 355 468
rect 355 467 356 468
rect 356 467 357 468
rect 357 467 358 468
rect 358 467 359 468
rect 359 467 360 468
rect 360 467 361 468
rect 361 467 362 468
rect 362 467 363 468
rect 363 467 364 468
rect 364 467 365 468
rect 365 467 366 468
rect 366 467 367 468
rect 367 467 368 468
rect 368 467 369 468
rect 369 467 370 468
rect 370 467 371 468
rect 371 467 372 468
rect 372 467 373 468
rect 373 467 374 468
rect 409 467 410 468
rect 410 467 411 468
rect 411 467 412 468
rect 412 467 413 468
rect 413 467 414 468
rect 414 467 415 468
rect 415 467 416 468
rect 416 467 417 468
rect 417 467 418 468
rect 418 467 419 468
rect 419 467 420 468
rect 420 467 421 468
rect 203 466 204 467
rect 204 466 205 467
rect 205 466 206 467
rect 206 466 207 467
rect 207 466 208 467
rect 208 466 209 467
rect 347 466 348 467
rect 348 466 349 467
rect 349 466 350 467
rect 350 466 351 467
rect 351 466 352 467
rect 352 466 353 467
rect 353 466 354 467
rect 354 466 355 467
rect 355 466 356 467
rect 356 466 357 467
rect 357 466 358 467
rect 358 466 359 467
rect 359 466 360 467
rect 360 466 361 467
rect 361 466 362 467
rect 362 466 363 467
rect 363 466 364 467
rect 364 466 365 467
rect 365 466 366 467
rect 366 466 367 467
rect 367 466 368 467
rect 368 466 369 467
rect 369 466 370 467
rect 370 466 371 467
rect 371 466 372 467
rect 372 466 373 467
rect 373 466 374 467
rect 407 466 408 467
rect 408 466 409 467
rect 409 466 410 467
rect 410 466 411 467
rect 411 466 412 467
rect 412 466 413 467
rect 413 466 414 467
rect 414 466 415 467
rect 415 466 416 467
rect 416 466 417 467
rect 417 466 418 467
rect 418 466 419 467
rect 419 466 420 467
rect 420 466 421 467
rect 203 465 204 466
rect 204 465 205 466
rect 205 465 206 466
rect 206 465 207 466
rect 347 465 348 466
rect 348 465 349 466
rect 349 465 350 466
rect 350 465 351 466
rect 351 465 352 466
rect 352 465 353 466
rect 353 465 354 466
rect 354 465 355 466
rect 355 465 356 466
rect 356 465 357 466
rect 357 465 358 466
rect 358 465 359 466
rect 359 465 360 466
rect 360 465 361 466
rect 361 465 362 466
rect 362 465 363 466
rect 363 465 364 466
rect 364 465 365 466
rect 365 465 366 466
rect 366 465 367 466
rect 367 465 368 466
rect 368 465 369 466
rect 369 465 370 466
rect 370 465 371 466
rect 371 465 372 466
rect 372 465 373 466
rect 373 465 374 466
rect 407 465 408 466
rect 408 465 409 466
rect 409 465 410 466
rect 410 465 411 466
rect 411 465 412 466
rect 412 465 413 466
rect 413 465 414 466
rect 414 465 415 466
rect 415 465 416 466
rect 416 465 417 466
rect 199 464 200 465
rect 200 464 201 465
rect 201 464 202 465
rect 202 464 203 465
rect 203 464 204 465
rect 204 464 205 465
rect 205 464 206 465
rect 206 464 207 465
rect 345 464 346 465
rect 346 464 347 465
rect 347 464 348 465
rect 348 464 349 465
rect 349 464 350 465
rect 350 464 351 465
rect 351 464 352 465
rect 352 464 353 465
rect 353 464 354 465
rect 354 464 355 465
rect 355 464 356 465
rect 356 464 357 465
rect 357 464 358 465
rect 358 464 359 465
rect 359 464 360 465
rect 360 464 361 465
rect 361 464 362 465
rect 362 464 363 465
rect 363 464 364 465
rect 364 464 365 465
rect 365 464 366 465
rect 366 464 367 465
rect 367 464 368 465
rect 368 464 369 465
rect 369 464 370 465
rect 370 464 371 465
rect 371 464 372 465
rect 372 464 373 465
rect 373 464 374 465
rect 407 464 408 465
rect 408 464 409 465
rect 409 464 410 465
rect 410 464 411 465
rect 411 464 412 465
rect 412 464 413 465
rect 413 464 414 465
rect 414 464 415 465
rect 415 464 416 465
rect 416 464 417 465
rect 199 463 200 464
rect 200 463 201 464
rect 201 463 202 464
rect 202 463 203 464
rect 203 463 204 464
rect 204 463 205 464
rect 205 463 206 464
rect 345 463 346 464
rect 346 463 347 464
rect 347 463 348 464
rect 348 463 349 464
rect 349 463 350 464
rect 350 463 351 464
rect 351 463 352 464
rect 352 463 353 464
rect 353 463 354 464
rect 354 463 355 464
rect 355 463 356 464
rect 356 463 357 464
rect 357 463 358 464
rect 358 463 359 464
rect 359 463 360 464
rect 360 463 361 464
rect 361 463 362 464
rect 362 463 363 464
rect 363 463 364 464
rect 364 463 365 464
rect 365 463 366 464
rect 366 463 367 464
rect 367 463 368 464
rect 368 463 369 464
rect 369 463 370 464
rect 370 463 371 464
rect 371 463 372 464
rect 407 463 408 464
rect 408 463 409 464
rect 409 463 410 464
rect 410 463 411 464
rect 411 463 412 464
rect 412 463 413 464
rect 413 463 414 464
rect 414 463 415 464
rect 199 462 200 463
rect 200 462 201 463
rect 201 462 202 463
rect 202 462 203 463
rect 203 462 204 463
rect 204 462 205 463
rect 205 462 206 463
rect 345 462 346 463
rect 346 462 347 463
rect 347 462 348 463
rect 348 462 349 463
rect 349 462 350 463
rect 350 462 351 463
rect 351 462 352 463
rect 352 462 353 463
rect 353 462 354 463
rect 354 462 355 463
rect 355 462 356 463
rect 356 462 357 463
rect 357 462 358 463
rect 358 462 359 463
rect 359 462 360 463
rect 360 462 361 463
rect 361 462 362 463
rect 362 462 363 463
rect 363 462 364 463
rect 364 462 365 463
rect 365 462 366 463
rect 366 462 367 463
rect 367 462 368 463
rect 368 462 369 463
rect 369 462 370 463
rect 370 462 371 463
rect 371 462 372 463
rect 403 462 404 463
rect 404 462 405 463
rect 405 462 406 463
rect 406 462 407 463
rect 407 462 408 463
rect 408 462 409 463
rect 409 462 410 463
rect 410 462 411 463
rect 411 462 412 463
rect 412 462 413 463
rect 413 462 414 463
rect 414 462 415 463
rect 199 461 200 462
rect 200 461 201 462
rect 201 461 202 462
rect 345 461 346 462
rect 346 461 347 462
rect 347 461 348 462
rect 348 461 349 462
rect 349 461 350 462
rect 350 461 351 462
rect 351 461 352 462
rect 352 461 353 462
rect 353 461 354 462
rect 354 461 355 462
rect 355 461 356 462
rect 356 461 357 462
rect 357 461 358 462
rect 358 461 359 462
rect 359 461 360 462
rect 360 461 361 462
rect 361 461 362 462
rect 362 461 363 462
rect 363 461 364 462
rect 364 461 365 462
rect 365 461 366 462
rect 366 461 367 462
rect 367 461 368 462
rect 368 461 369 462
rect 369 461 370 462
rect 403 461 404 462
rect 404 461 405 462
rect 405 461 406 462
rect 406 461 407 462
rect 407 461 408 462
rect 408 461 409 462
rect 409 461 410 462
rect 410 461 411 462
rect 411 461 412 462
rect 195 460 196 461
rect 196 460 197 461
rect 197 460 198 461
rect 198 460 199 461
rect 199 460 200 461
rect 200 460 201 461
rect 201 460 202 461
rect 345 460 346 461
rect 346 460 347 461
rect 347 460 348 461
rect 348 460 349 461
rect 349 460 350 461
rect 350 460 351 461
rect 351 460 352 461
rect 352 460 353 461
rect 353 460 354 461
rect 354 460 355 461
rect 355 460 356 461
rect 356 460 357 461
rect 357 460 358 461
rect 358 460 359 461
rect 359 460 360 461
rect 360 460 361 461
rect 361 460 362 461
rect 362 460 363 461
rect 363 460 364 461
rect 364 460 365 461
rect 365 460 366 461
rect 366 460 367 461
rect 367 460 368 461
rect 368 460 369 461
rect 369 460 370 461
rect 401 460 402 461
rect 402 460 403 461
rect 403 460 404 461
rect 404 460 405 461
rect 405 460 406 461
rect 406 460 407 461
rect 407 460 408 461
rect 408 460 409 461
rect 409 460 410 461
rect 410 460 411 461
rect 411 460 412 461
rect 195 459 196 460
rect 196 459 197 460
rect 197 459 198 460
rect 198 459 199 460
rect 199 459 200 460
rect 200 459 201 460
rect 201 459 202 460
rect 345 459 346 460
rect 346 459 347 460
rect 347 459 348 460
rect 348 459 349 460
rect 349 459 350 460
rect 350 459 351 460
rect 351 459 352 460
rect 352 459 353 460
rect 353 459 354 460
rect 354 459 355 460
rect 355 459 356 460
rect 356 459 357 460
rect 357 459 358 460
rect 358 459 359 460
rect 359 459 360 460
rect 360 459 361 460
rect 361 459 362 460
rect 362 459 363 460
rect 363 459 364 460
rect 364 459 365 460
rect 365 459 366 460
rect 366 459 367 460
rect 367 459 368 460
rect 368 459 369 460
rect 369 459 370 460
rect 401 459 402 460
rect 402 459 403 460
rect 403 459 404 460
rect 404 459 405 460
rect 405 459 406 460
rect 406 459 407 460
rect 407 459 408 460
rect 408 459 409 460
rect 409 459 410 460
rect 193 458 194 459
rect 194 458 195 459
rect 195 458 196 459
rect 196 458 197 459
rect 197 458 198 459
rect 198 458 199 459
rect 199 458 200 459
rect 200 458 201 459
rect 201 458 202 459
rect 343 458 344 459
rect 344 458 345 459
rect 345 458 346 459
rect 346 458 347 459
rect 347 458 348 459
rect 348 458 349 459
rect 349 458 350 459
rect 350 458 351 459
rect 351 458 352 459
rect 352 458 353 459
rect 353 458 354 459
rect 354 458 355 459
rect 355 458 356 459
rect 356 458 357 459
rect 357 458 358 459
rect 358 458 359 459
rect 359 458 360 459
rect 360 458 361 459
rect 361 458 362 459
rect 362 458 363 459
rect 363 458 364 459
rect 364 458 365 459
rect 365 458 366 459
rect 366 458 367 459
rect 367 458 368 459
rect 368 458 369 459
rect 369 458 370 459
rect 399 458 400 459
rect 400 458 401 459
rect 401 458 402 459
rect 402 458 403 459
rect 403 458 404 459
rect 404 458 405 459
rect 405 458 406 459
rect 406 458 407 459
rect 407 458 408 459
rect 408 458 409 459
rect 409 458 410 459
rect 193 457 194 458
rect 194 457 195 458
rect 195 457 196 458
rect 196 457 197 458
rect 197 457 198 458
rect 343 457 344 458
rect 344 457 345 458
rect 345 457 346 458
rect 346 457 347 458
rect 347 457 348 458
rect 348 457 349 458
rect 349 457 350 458
rect 350 457 351 458
rect 351 457 352 458
rect 352 457 353 458
rect 353 457 354 458
rect 354 457 355 458
rect 355 457 356 458
rect 356 457 357 458
rect 357 457 358 458
rect 358 457 359 458
rect 359 457 360 458
rect 360 457 361 458
rect 361 457 362 458
rect 362 457 363 458
rect 363 457 364 458
rect 364 457 365 458
rect 365 457 366 458
rect 366 457 367 458
rect 367 457 368 458
rect 368 457 369 458
rect 399 457 400 458
rect 400 457 401 458
rect 401 457 402 458
rect 402 457 403 458
rect 403 457 404 458
rect 404 457 405 458
rect 405 457 406 458
rect 193 456 194 457
rect 194 456 195 457
rect 195 456 196 457
rect 196 456 197 457
rect 197 456 198 457
rect 343 456 344 457
rect 344 456 345 457
rect 345 456 346 457
rect 346 456 347 457
rect 347 456 348 457
rect 348 456 349 457
rect 349 456 350 457
rect 350 456 351 457
rect 351 456 352 457
rect 352 456 353 457
rect 353 456 354 457
rect 354 456 355 457
rect 355 456 356 457
rect 356 456 357 457
rect 357 456 358 457
rect 358 456 359 457
rect 359 456 360 457
rect 360 456 361 457
rect 361 456 362 457
rect 362 456 363 457
rect 363 456 364 457
rect 364 456 365 457
rect 365 456 366 457
rect 366 456 367 457
rect 367 456 368 457
rect 368 456 369 457
rect 397 456 398 457
rect 398 456 399 457
rect 399 456 400 457
rect 400 456 401 457
rect 401 456 402 457
rect 402 456 403 457
rect 403 456 404 457
rect 404 456 405 457
rect 405 456 406 457
rect 193 455 194 456
rect 194 455 195 456
rect 195 455 196 456
rect 343 455 344 456
rect 344 455 345 456
rect 345 455 346 456
rect 346 455 347 456
rect 347 455 348 456
rect 348 455 349 456
rect 349 455 350 456
rect 350 455 351 456
rect 351 455 352 456
rect 352 455 353 456
rect 353 455 354 456
rect 354 455 355 456
rect 355 455 356 456
rect 356 455 357 456
rect 357 455 358 456
rect 358 455 359 456
rect 359 455 360 456
rect 360 455 361 456
rect 361 455 362 456
rect 362 455 363 456
rect 363 455 364 456
rect 364 455 365 456
rect 365 455 366 456
rect 366 455 367 456
rect 397 455 398 456
rect 398 455 399 456
rect 399 455 400 456
rect 400 455 401 456
rect 401 455 402 456
rect 402 455 403 456
rect 403 455 404 456
rect 190 454 191 455
rect 191 454 192 455
rect 192 454 193 455
rect 193 454 194 455
rect 194 454 195 455
rect 195 454 196 455
rect 343 454 344 455
rect 344 454 345 455
rect 345 454 346 455
rect 346 454 347 455
rect 347 454 348 455
rect 348 454 349 455
rect 349 454 350 455
rect 350 454 351 455
rect 351 454 352 455
rect 352 454 353 455
rect 353 454 354 455
rect 354 454 355 455
rect 355 454 356 455
rect 356 454 357 455
rect 357 454 358 455
rect 358 454 359 455
rect 359 454 360 455
rect 360 454 361 455
rect 361 454 362 455
rect 362 454 363 455
rect 363 454 364 455
rect 364 454 365 455
rect 365 454 366 455
rect 366 454 367 455
rect 394 454 395 455
rect 395 454 396 455
rect 396 454 397 455
rect 397 454 398 455
rect 398 454 399 455
rect 399 454 400 455
rect 400 454 401 455
rect 401 454 402 455
rect 402 454 403 455
rect 403 454 404 455
rect 190 453 191 454
rect 191 453 192 454
rect 192 453 193 454
rect 193 453 194 454
rect 343 453 344 454
rect 344 453 345 454
rect 345 453 346 454
rect 346 453 347 454
rect 347 453 348 454
rect 348 453 349 454
rect 349 453 350 454
rect 350 453 351 454
rect 351 453 352 454
rect 352 453 353 454
rect 353 453 354 454
rect 354 453 355 454
rect 355 453 356 454
rect 356 453 357 454
rect 357 453 358 454
rect 358 453 359 454
rect 359 453 360 454
rect 360 453 361 454
rect 361 453 362 454
rect 362 453 363 454
rect 363 453 364 454
rect 364 453 365 454
rect 365 453 366 454
rect 366 453 367 454
rect 394 453 395 454
rect 395 453 396 454
rect 396 453 397 454
rect 397 453 398 454
rect 398 453 399 454
rect 399 453 400 454
rect 400 453 401 454
rect 401 453 402 454
rect 188 452 189 453
rect 189 452 190 453
rect 190 452 191 453
rect 191 452 192 453
rect 192 452 193 453
rect 193 452 194 453
rect 341 452 342 453
rect 342 452 343 453
rect 343 452 344 453
rect 344 452 345 453
rect 345 452 346 453
rect 346 452 347 453
rect 347 452 348 453
rect 348 452 349 453
rect 349 452 350 453
rect 350 452 351 453
rect 351 452 352 453
rect 352 452 353 453
rect 353 452 354 453
rect 354 452 355 453
rect 355 452 356 453
rect 356 452 357 453
rect 357 452 358 453
rect 358 452 359 453
rect 359 452 360 453
rect 360 452 361 453
rect 361 452 362 453
rect 362 452 363 453
rect 363 452 364 453
rect 364 452 365 453
rect 365 452 366 453
rect 366 452 367 453
rect 392 452 393 453
rect 393 452 394 453
rect 394 452 395 453
rect 395 452 396 453
rect 396 452 397 453
rect 397 452 398 453
rect 398 452 399 453
rect 399 452 400 453
rect 400 452 401 453
rect 401 452 402 453
rect 188 451 189 452
rect 189 451 190 452
rect 190 451 191 452
rect 191 451 192 452
rect 192 451 193 452
rect 193 451 194 452
rect 341 451 342 452
rect 342 451 343 452
rect 343 451 344 452
rect 344 451 345 452
rect 345 451 346 452
rect 346 451 347 452
rect 347 451 348 452
rect 348 451 349 452
rect 349 451 350 452
rect 350 451 351 452
rect 351 451 352 452
rect 352 451 353 452
rect 353 451 354 452
rect 354 451 355 452
rect 355 451 356 452
rect 356 451 357 452
rect 357 451 358 452
rect 358 451 359 452
rect 359 451 360 452
rect 360 451 361 452
rect 361 451 362 452
rect 362 451 363 452
rect 363 451 364 452
rect 364 451 365 452
rect 392 451 393 452
rect 393 451 394 452
rect 394 451 395 452
rect 395 451 396 452
rect 396 451 397 452
rect 397 451 398 452
rect 186 450 187 451
rect 187 450 188 451
rect 188 450 189 451
rect 189 450 190 451
rect 190 450 191 451
rect 191 450 192 451
rect 192 450 193 451
rect 193 450 194 451
rect 341 450 342 451
rect 342 450 343 451
rect 343 450 344 451
rect 344 450 345 451
rect 345 450 346 451
rect 346 450 347 451
rect 347 450 348 451
rect 348 450 349 451
rect 349 450 350 451
rect 350 450 351 451
rect 351 450 352 451
rect 352 450 353 451
rect 353 450 354 451
rect 354 450 355 451
rect 355 450 356 451
rect 356 450 357 451
rect 357 450 358 451
rect 358 450 359 451
rect 359 450 360 451
rect 360 450 361 451
rect 361 450 362 451
rect 362 450 363 451
rect 363 450 364 451
rect 364 450 365 451
rect 390 450 391 451
rect 391 450 392 451
rect 392 450 393 451
rect 393 450 394 451
rect 394 450 395 451
rect 395 450 396 451
rect 396 450 397 451
rect 397 450 398 451
rect 186 449 187 450
rect 187 449 188 450
rect 188 449 189 450
rect 189 449 190 450
rect 190 449 191 450
rect 341 449 342 450
rect 342 449 343 450
rect 343 449 344 450
rect 344 449 345 450
rect 345 449 346 450
rect 346 449 347 450
rect 347 449 348 450
rect 348 449 349 450
rect 349 449 350 450
rect 350 449 351 450
rect 351 449 352 450
rect 352 449 353 450
rect 353 449 354 450
rect 354 449 355 450
rect 355 449 356 450
rect 356 449 357 450
rect 357 449 358 450
rect 358 449 359 450
rect 359 449 360 450
rect 360 449 361 450
rect 361 449 362 450
rect 362 449 363 450
rect 390 449 391 450
rect 391 449 392 450
rect 392 449 393 450
rect 393 449 394 450
rect 394 449 395 450
rect 395 449 396 450
rect 396 449 397 450
rect 397 449 398 450
rect 184 448 185 449
rect 185 448 186 449
rect 186 448 187 449
rect 187 448 188 449
rect 188 448 189 449
rect 189 448 190 449
rect 190 448 191 449
rect 341 448 342 449
rect 342 448 343 449
rect 343 448 344 449
rect 344 448 345 449
rect 345 448 346 449
rect 346 448 347 449
rect 347 448 348 449
rect 348 448 349 449
rect 349 448 350 449
rect 350 448 351 449
rect 351 448 352 449
rect 352 448 353 449
rect 353 448 354 449
rect 354 448 355 449
rect 355 448 356 449
rect 356 448 357 449
rect 357 448 358 449
rect 358 448 359 449
rect 359 448 360 449
rect 360 448 361 449
rect 361 448 362 449
rect 362 448 363 449
rect 386 448 387 449
rect 387 448 388 449
rect 388 448 389 449
rect 389 448 390 449
rect 390 448 391 449
rect 391 448 392 449
rect 392 448 393 449
rect 393 448 394 449
rect 394 448 395 449
rect 395 448 396 449
rect 396 448 397 449
rect 397 448 398 449
rect 184 447 185 448
rect 185 447 186 448
rect 186 447 187 448
rect 187 447 188 448
rect 188 447 189 448
rect 341 447 342 448
rect 342 447 343 448
rect 343 447 344 448
rect 344 447 345 448
rect 345 447 346 448
rect 346 447 347 448
rect 347 447 348 448
rect 348 447 349 448
rect 349 447 350 448
rect 350 447 351 448
rect 351 447 352 448
rect 352 447 353 448
rect 353 447 354 448
rect 354 447 355 448
rect 355 447 356 448
rect 356 447 357 448
rect 357 447 358 448
rect 358 447 359 448
rect 359 447 360 448
rect 360 447 361 448
rect 361 447 362 448
rect 362 447 363 448
rect 386 447 387 448
rect 387 447 388 448
rect 388 447 389 448
rect 389 447 390 448
rect 390 447 391 448
rect 391 447 392 448
rect 392 447 393 448
rect 393 447 394 448
rect 394 447 395 448
rect 182 446 183 447
rect 183 446 184 447
rect 184 446 185 447
rect 185 446 186 447
rect 186 446 187 447
rect 187 446 188 447
rect 188 446 189 447
rect 341 446 342 447
rect 342 446 343 447
rect 343 446 344 447
rect 344 446 345 447
rect 345 446 346 447
rect 346 446 347 447
rect 347 446 348 447
rect 348 446 349 447
rect 349 446 350 447
rect 350 446 351 447
rect 351 446 352 447
rect 352 446 353 447
rect 353 446 354 447
rect 354 446 355 447
rect 355 446 356 447
rect 356 446 357 447
rect 357 446 358 447
rect 358 446 359 447
rect 359 446 360 447
rect 360 446 361 447
rect 361 446 362 447
rect 362 446 363 447
rect 384 446 385 447
rect 385 446 386 447
rect 386 446 387 447
rect 387 446 388 447
rect 388 446 389 447
rect 389 446 390 447
rect 390 446 391 447
rect 391 446 392 447
rect 392 446 393 447
rect 393 446 394 447
rect 394 446 395 447
rect 182 445 183 446
rect 183 445 184 446
rect 184 445 185 446
rect 185 445 186 446
rect 186 445 187 446
rect 341 445 342 446
rect 342 445 343 446
rect 343 445 344 446
rect 344 445 345 446
rect 345 445 346 446
rect 346 445 347 446
rect 347 445 348 446
rect 348 445 349 446
rect 349 445 350 446
rect 350 445 351 446
rect 351 445 352 446
rect 352 445 353 446
rect 353 445 354 446
rect 354 445 355 446
rect 355 445 356 446
rect 356 445 357 446
rect 357 445 358 446
rect 358 445 359 446
rect 359 445 360 446
rect 360 445 361 446
rect 384 445 385 446
rect 385 445 386 446
rect 386 445 387 446
rect 387 445 388 446
rect 388 445 389 446
rect 389 445 390 446
rect 390 445 391 446
rect 391 445 392 446
rect 392 445 393 446
rect 180 444 181 445
rect 181 444 182 445
rect 182 444 183 445
rect 183 444 184 445
rect 184 444 185 445
rect 185 444 186 445
rect 186 444 187 445
rect 341 444 342 445
rect 342 444 343 445
rect 343 444 344 445
rect 344 444 345 445
rect 345 444 346 445
rect 346 444 347 445
rect 347 444 348 445
rect 348 444 349 445
rect 349 444 350 445
rect 350 444 351 445
rect 351 444 352 445
rect 352 444 353 445
rect 353 444 354 445
rect 354 444 355 445
rect 355 444 356 445
rect 356 444 357 445
rect 357 444 358 445
rect 358 444 359 445
rect 359 444 360 445
rect 360 444 361 445
rect 381 444 382 445
rect 382 444 383 445
rect 383 444 384 445
rect 384 444 385 445
rect 385 444 386 445
rect 386 444 387 445
rect 387 444 388 445
rect 388 444 389 445
rect 389 444 390 445
rect 390 444 391 445
rect 391 444 392 445
rect 392 444 393 445
rect 180 443 181 444
rect 181 443 182 444
rect 182 443 183 444
rect 183 443 184 444
rect 184 443 185 444
rect 341 443 342 444
rect 342 443 343 444
rect 343 443 344 444
rect 344 443 345 444
rect 345 443 346 444
rect 346 443 347 444
rect 347 443 348 444
rect 348 443 349 444
rect 349 443 350 444
rect 350 443 351 444
rect 351 443 352 444
rect 352 443 353 444
rect 353 443 354 444
rect 354 443 355 444
rect 355 443 356 444
rect 356 443 357 444
rect 357 443 358 444
rect 358 443 359 444
rect 359 443 360 444
rect 360 443 361 444
rect 381 443 382 444
rect 382 443 383 444
rect 383 443 384 444
rect 384 443 385 444
rect 385 443 386 444
rect 386 443 387 444
rect 387 443 388 444
rect 388 443 389 444
rect 389 443 390 444
rect 390 443 391 444
rect 178 442 179 443
rect 179 442 180 443
rect 180 442 181 443
rect 181 442 182 443
rect 182 442 183 443
rect 183 442 184 443
rect 184 442 185 443
rect 341 442 342 443
rect 342 442 343 443
rect 343 442 344 443
rect 344 442 345 443
rect 345 442 346 443
rect 346 442 347 443
rect 347 442 348 443
rect 348 442 349 443
rect 349 442 350 443
rect 350 442 351 443
rect 351 442 352 443
rect 352 442 353 443
rect 353 442 354 443
rect 354 442 355 443
rect 355 442 356 443
rect 356 442 357 443
rect 357 442 358 443
rect 358 442 359 443
rect 359 442 360 443
rect 360 442 361 443
rect 379 442 380 443
rect 380 442 381 443
rect 381 442 382 443
rect 382 442 383 443
rect 383 442 384 443
rect 384 442 385 443
rect 385 442 386 443
rect 386 442 387 443
rect 387 442 388 443
rect 388 442 389 443
rect 389 442 390 443
rect 390 442 391 443
rect 178 441 179 442
rect 179 441 180 442
rect 180 441 181 442
rect 181 441 182 442
rect 182 441 183 442
rect 341 441 342 442
rect 342 441 343 442
rect 343 441 344 442
rect 344 441 345 442
rect 345 441 346 442
rect 346 441 347 442
rect 347 441 348 442
rect 348 441 349 442
rect 349 441 350 442
rect 350 441 351 442
rect 351 441 352 442
rect 352 441 353 442
rect 353 441 354 442
rect 354 441 355 442
rect 355 441 356 442
rect 356 441 357 442
rect 357 441 358 442
rect 358 441 359 442
rect 379 441 380 442
rect 380 441 381 442
rect 381 441 382 442
rect 382 441 383 442
rect 383 441 384 442
rect 384 441 385 442
rect 385 441 386 442
rect 386 441 387 442
rect 387 441 388 442
rect 388 441 389 442
rect 175 440 176 441
rect 176 440 177 441
rect 177 440 178 441
rect 178 440 179 441
rect 179 440 180 441
rect 180 440 181 441
rect 181 440 182 441
rect 182 440 183 441
rect 339 440 340 441
rect 340 440 341 441
rect 341 440 342 441
rect 342 440 343 441
rect 343 440 344 441
rect 344 440 345 441
rect 345 440 346 441
rect 346 440 347 441
rect 347 440 348 441
rect 348 440 349 441
rect 349 440 350 441
rect 350 440 351 441
rect 351 440 352 441
rect 352 440 353 441
rect 353 440 354 441
rect 354 440 355 441
rect 355 440 356 441
rect 356 440 357 441
rect 357 440 358 441
rect 358 440 359 441
rect 375 440 376 441
rect 376 440 377 441
rect 377 440 378 441
rect 378 440 379 441
rect 379 440 380 441
rect 380 440 381 441
rect 381 440 382 441
rect 382 440 383 441
rect 383 440 384 441
rect 384 440 385 441
rect 385 440 386 441
rect 386 440 387 441
rect 387 440 388 441
rect 388 440 389 441
rect 175 439 176 440
rect 176 439 177 440
rect 177 439 178 440
rect 178 439 179 440
rect 339 439 340 440
rect 340 439 341 440
rect 341 439 342 440
rect 342 439 343 440
rect 343 439 344 440
rect 344 439 345 440
rect 345 439 346 440
rect 346 439 347 440
rect 347 439 348 440
rect 348 439 349 440
rect 349 439 350 440
rect 350 439 351 440
rect 351 439 352 440
rect 352 439 353 440
rect 353 439 354 440
rect 354 439 355 440
rect 355 439 356 440
rect 356 439 357 440
rect 357 439 358 440
rect 358 439 359 440
rect 375 439 376 440
rect 376 439 377 440
rect 377 439 378 440
rect 378 439 379 440
rect 379 439 380 440
rect 380 439 381 440
rect 381 439 382 440
rect 382 439 383 440
rect 383 439 384 440
rect 384 439 385 440
rect 385 439 386 440
rect 386 439 387 440
rect 173 438 174 439
rect 174 438 175 439
rect 175 438 176 439
rect 176 438 177 439
rect 177 438 178 439
rect 178 438 179 439
rect 339 438 340 439
rect 340 438 341 439
rect 341 438 342 439
rect 342 438 343 439
rect 343 438 344 439
rect 344 438 345 439
rect 345 438 346 439
rect 346 438 347 439
rect 347 438 348 439
rect 348 438 349 439
rect 349 438 350 439
rect 350 438 351 439
rect 351 438 352 439
rect 352 438 353 439
rect 353 438 354 439
rect 354 438 355 439
rect 355 438 356 439
rect 356 438 357 439
rect 357 438 358 439
rect 358 438 359 439
rect 373 438 374 439
rect 374 438 375 439
rect 375 438 376 439
rect 376 438 377 439
rect 377 438 378 439
rect 378 438 379 439
rect 379 438 380 439
rect 380 438 381 439
rect 381 438 382 439
rect 382 438 383 439
rect 383 438 384 439
rect 384 438 385 439
rect 385 438 386 439
rect 386 438 387 439
rect 173 437 174 438
rect 174 437 175 438
rect 175 437 176 438
rect 176 437 177 438
rect 341 437 342 438
rect 342 437 343 438
rect 343 437 344 438
rect 344 437 345 438
rect 345 437 346 438
rect 346 437 347 438
rect 347 437 348 438
rect 348 437 349 438
rect 349 437 350 438
rect 350 437 351 438
rect 351 437 352 438
rect 352 437 353 438
rect 353 437 354 438
rect 354 437 355 438
rect 355 437 356 438
rect 356 437 357 438
rect 357 437 358 438
rect 358 437 359 438
rect 373 437 374 438
rect 374 437 375 438
rect 375 437 376 438
rect 376 437 377 438
rect 377 437 378 438
rect 378 437 379 438
rect 379 437 380 438
rect 380 437 381 438
rect 381 437 382 438
rect 382 437 383 438
rect 383 437 384 438
rect 384 437 385 438
rect 385 437 386 438
rect 386 437 387 438
rect 171 436 172 437
rect 172 436 173 437
rect 173 436 174 437
rect 174 436 175 437
rect 175 436 176 437
rect 176 436 177 437
rect 341 436 342 437
rect 342 436 343 437
rect 343 436 344 437
rect 344 436 345 437
rect 345 436 346 437
rect 346 436 347 437
rect 347 436 348 437
rect 348 436 349 437
rect 349 436 350 437
rect 350 436 351 437
rect 351 436 352 437
rect 352 436 353 437
rect 353 436 354 437
rect 354 436 355 437
rect 355 436 356 437
rect 356 436 357 437
rect 357 436 358 437
rect 358 436 359 437
rect 371 436 372 437
rect 372 436 373 437
rect 373 436 374 437
rect 374 436 375 437
rect 375 436 376 437
rect 376 436 377 437
rect 377 436 378 437
rect 378 436 379 437
rect 379 436 380 437
rect 380 436 381 437
rect 381 436 382 437
rect 382 436 383 437
rect 383 436 384 437
rect 384 436 385 437
rect 385 436 386 437
rect 386 436 387 437
rect 171 435 172 436
rect 172 435 173 436
rect 173 435 174 436
rect 174 435 175 436
rect 175 435 176 436
rect 341 435 342 436
rect 342 435 343 436
rect 343 435 344 436
rect 344 435 345 436
rect 345 435 346 436
rect 346 435 347 436
rect 347 435 348 436
rect 348 435 349 436
rect 349 435 350 436
rect 350 435 351 436
rect 351 435 352 436
rect 352 435 353 436
rect 353 435 354 436
rect 354 435 355 436
rect 355 435 356 436
rect 356 435 357 436
rect 371 435 372 436
rect 372 435 373 436
rect 373 435 374 436
rect 374 435 375 436
rect 375 435 376 436
rect 376 435 377 436
rect 377 435 378 436
rect 378 435 379 436
rect 379 435 380 436
rect 380 435 381 436
rect 381 435 382 436
rect 382 435 383 436
rect 383 435 384 436
rect 384 435 385 436
rect 169 434 170 435
rect 170 434 171 435
rect 171 434 172 435
rect 172 434 173 435
rect 173 434 174 435
rect 174 434 175 435
rect 175 434 176 435
rect 341 434 342 435
rect 342 434 343 435
rect 343 434 344 435
rect 344 434 345 435
rect 345 434 346 435
rect 346 434 347 435
rect 347 434 348 435
rect 348 434 349 435
rect 349 434 350 435
rect 350 434 351 435
rect 351 434 352 435
rect 352 434 353 435
rect 353 434 354 435
rect 354 434 355 435
rect 355 434 356 435
rect 356 434 357 435
rect 369 434 370 435
rect 370 434 371 435
rect 371 434 372 435
rect 372 434 373 435
rect 373 434 374 435
rect 374 434 375 435
rect 375 434 376 435
rect 376 434 377 435
rect 377 434 378 435
rect 378 434 379 435
rect 379 434 380 435
rect 380 434 381 435
rect 381 434 382 435
rect 382 434 383 435
rect 383 434 384 435
rect 384 434 385 435
rect 169 433 170 434
rect 170 433 171 434
rect 171 433 172 434
rect 341 433 342 434
rect 342 433 343 434
rect 343 433 344 434
rect 344 433 345 434
rect 345 433 346 434
rect 346 433 347 434
rect 347 433 348 434
rect 348 433 349 434
rect 349 433 350 434
rect 350 433 351 434
rect 351 433 352 434
rect 352 433 353 434
rect 353 433 354 434
rect 354 433 355 434
rect 355 433 356 434
rect 356 433 357 434
rect 369 433 370 434
rect 370 433 371 434
rect 371 433 372 434
rect 372 433 373 434
rect 373 433 374 434
rect 374 433 375 434
rect 375 433 376 434
rect 376 433 377 434
rect 377 433 378 434
rect 378 433 379 434
rect 379 433 380 434
rect 380 433 381 434
rect 381 433 382 434
rect 382 433 383 434
rect 383 433 384 434
rect 169 432 170 433
rect 170 432 171 433
rect 171 432 172 433
rect 341 432 342 433
rect 342 432 343 433
rect 343 432 344 433
rect 344 432 345 433
rect 345 432 346 433
rect 346 432 347 433
rect 347 432 348 433
rect 348 432 349 433
rect 349 432 350 433
rect 350 432 351 433
rect 351 432 352 433
rect 352 432 353 433
rect 353 432 354 433
rect 354 432 355 433
rect 355 432 356 433
rect 356 432 357 433
rect 369 432 370 433
rect 370 432 371 433
rect 371 432 372 433
rect 372 432 373 433
rect 373 432 374 433
rect 374 432 375 433
rect 375 432 376 433
rect 376 432 377 433
rect 377 432 378 433
rect 378 432 379 433
rect 379 432 380 433
rect 380 432 381 433
rect 381 432 382 433
rect 382 432 383 433
rect 383 432 384 433
rect 167 431 168 432
rect 168 431 169 432
rect 169 431 170 432
rect 170 431 171 432
rect 171 431 172 432
rect 341 431 342 432
rect 342 431 343 432
rect 343 431 344 432
rect 344 431 345 432
rect 345 431 346 432
rect 346 431 347 432
rect 347 431 348 432
rect 348 431 349 432
rect 349 431 350 432
rect 350 431 351 432
rect 351 431 352 432
rect 352 431 353 432
rect 353 431 354 432
rect 354 431 355 432
rect 355 431 356 432
rect 356 431 357 432
rect 368 431 369 432
rect 369 431 370 432
rect 370 431 371 432
rect 371 431 372 432
rect 372 431 373 432
rect 373 431 374 432
rect 374 431 375 432
rect 375 431 376 432
rect 376 431 377 432
rect 377 431 378 432
rect 378 431 379 432
rect 379 431 380 432
rect 380 431 381 432
rect 381 431 382 432
rect 382 431 383 432
rect 383 431 384 432
rect 167 430 168 431
rect 168 430 169 431
rect 169 430 170 431
rect 341 430 342 431
rect 342 430 343 431
rect 343 430 344 431
rect 344 430 345 431
rect 345 430 346 431
rect 346 430 347 431
rect 347 430 348 431
rect 348 430 349 431
rect 349 430 350 431
rect 350 430 351 431
rect 351 430 352 431
rect 352 430 353 431
rect 353 430 354 431
rect 354 430 355 431
rect 368 430 369 431
rect 369 430 370 431
rect 370 430 371 431
rect 371 430 372 431
rect 372 430 373 431
rect 373 430 374 431
rect 374 430 375 431
rect 375 430 376 431
rect 376 430 377 431
rect 377 430 378 431
rect 378 430 379 431
rect 379 430 380 431
rect 380 430 381 431
rect 381 430 382 431
rect 165 429 166 430
rect 166 429 167 430
rect 167 429 168 430
rect 168 429 169 430
rect 169 429 170 430
rect 339 429 340 430
rect 340 429 341 430
rect 341 429 342 430
rect 342 429 343 430
rect 343 429 344 430
rect 344 429 345 430
rect 345 429 346 430
rect 346 429 347 430
rect 347 429 348 430
rect 348 429 349 430
rect 349 429 350 430
rect 350 429 351 430
rect 351 429 352 430
rect 352 429 353 430
rect 353 429 354 430
rect 354 429 355 430
rect 366 429 367 430
rect 367 429 368 430
rect 368 429 369 430
rect 369 429 370 430
rect 370 429 371 430
rect 371 429 372 430
rect 372 429 373 430
rect 373 429 374 430
rect 374 429 375 430
rect 375 429 376 430
rect 376 429 377 430
rect 377 429 378 430
rect 378 429 379 430
rect 379 429 380 430
rect 380 429 381 430
rect 381 429 382 430
rect 165 428 166 429
rect 166 428 167 429
rect 167 428 168 429
rect 339 428 340 429
rect 340 428 341 429
rect 341 428 342 429
rect 342 428 343 429
rect 343 428 344 429
rect 344 428 345 429
rect 345 428 346 429
rect 346 428 347 429
rect 347 428 348 429
rect 348 428 349 429
rect 349 428 350 429
rect 350 428 351 429
rect 351 428 352 429
rect 352 428 353 429
rect 353 428 354 429
rect 354 428 355 429
rect 366 428 367 429
rect 367 428 368 429
rect 368 428 369 429
rect 369 428 370 429
rect 370 428 371 429
rect 371 428 372 429
rect 372 428 373 429
rect 373 428 374 429
rect 374 428 375 429
rect 375 428 376 429
rect 376 428 377 429
rect 377 428 378 429
rect 378 428 379 429
rect 379 428 380 429
rect 162 427 163 428
rect 163 427 164 428
rect 164 427 165 428
rect 165 427 166 428
rect 166 427 167 428
rect 167 427 168 428
rect 339 427 340 428
rect 340 427 341 428
rect 341 427 342 428
rect 342 427 343 428
rect 343 427 344 428
rect 344 427 345 428
rect 345 427 346 428
rect 346 427 347 428
rect 347 427 348 428
rect 348 427 349 428
rect 349 427 350 428
rect 350 427 351 428
rect 351 427 352 428
rect 352 427 353 428
rect 353 427 354 428
rect 354 427 355 428
rect 364 427 365 428
rect 365 427 366 428
rect 366 427 367 428
rect 367 427 368 428
rect 368 427 369 428
rect 369 427 370 428
rect 370 427 371 428
rect 371 427 372 428
rect 372 427 373 428
rect 373 427 374 428
rect 374 427 375 428
rect 375 427 376 428
rect 376 427 377 428
rect 377 427 378 428
rect 378 427 379 428
rect 379 427 380 428
rect 162 426 163 427
rect 163 426 164 427
rect 164 426 165 427
rect 165 426 166 427
rect 339 426 340 427
rect 340 426 341 427
rect 341 426 342 427
rect 342 426 343 427
rect 343 426 344 427
rect 344 426 345 427
rect 345 426 346 427
rect 346 426 347 427
rect 347 426 348 427
rect 348 426 349 427
rect 349 426 350 427
rect 350 426 351 427
rect 351 426 352 427
rect 352 426 353 427
rect 353 426 354 427
rect 354 426 355 427
rect 364 426 365 427
rect 365 426 366 427
rect 366 426 367 427
rect 367 426 368 427
rect 368 426 369 427
rect 369 426 370 427
rect 370 426 371 427
rect 371 426 372 427
rect 372 426 373 427
rect 373 426 374 427
rect 374 426 375 427
rect 375 426 376 427
rect 376 426 377 427
rect 377 426 378 427
rect 160 425 161 426
rect 161 425 162 426
rect 162 425 163 426
rect 163 425 164 426
rect 164 425 165 426
rect 165 425 166 426
rect 235 425 236 426
rect 236 425 237 426
rect 242 425 243 426
rect 243 425 244 426
rect 244 425 245 426
rect 339 425 340 426
rect 340 425 341 426
rect 341 425 342 426
rect 342 425 343 426
rect 343 425 344 426
rect 344 425 345 426
rect 345 425 346 426
rect 346 425 347 426
rect 347 425 348 426
rect 348 425 349 426
rect 349 425 350 426
rect 350 425 351 426
rect 351 425 352 426
rect 352 425 353 426
rect 353 425 354 426
rect 354 425 355 426
rect 362 425 363 426
rect 363 425 364 426
rect 364 425 365 426
rect 365 425 366 426
rect 366 425 367 426
rect 367 425 368 426
rect 368 425 369 426
rect 369 425 370 426
rect 370 425 371 426
rect 371 425 372 426
rect 372 425 373 426
rect 373 425 374 426
rect 374 425 375 426
rect 375 425 376 426
rect 376 425 377 426
rect 377 425 378 426
rect 160 424 161 425
rect 161 424 162 425
rect 162 424 163 425
rect 235 424 236 425
rect 236 424 237 425
rect 242 424 243 425
rect 243 424 244 425
rect 244 424 245 425
rect 341 424 342 425
rect 342 424 343 425
rect 343 424 344 425
rect 344 424 345 425
rect 345 424 346 425
rect 346 424 347 425
rect 347 424 348 425
rect 348 424 349 425
rect 349 424 350 425
rect 350 424 351 425
rect 351 424 352 425
rect 352 424 353 425
rect 353 424 354 425
rect 362 424 363 425
rect 363 424 364 425
rect 364 424 365 425
rect 365 424 366 425
rect 366 424 367 425
rect 367 424 368 425
rect 368 424 369 425
rect 369 424 370 425
rect 370 424 371 425
rect 371 424 372 425
rect 372 424 373 425
rect 373 424 374 425
rect 374 424 375 425
rect 375 424 376 425
rect 376 424 377 425
rect 377 424 378 425
rect 158 423 159 424
rect 159 423 160 424
rect 160 423 161 424
rect 161 423 162 424
rect 162 423 163 424
rect 221 423 222 424
rect 222 423 223 424
rect 223 423 224 424
rect 224 423 225 424
rect 225 423 226 424
rect 226 423 227 424
rect 227 423 228 424
rect 228 423 229 424
rect 229 423 230 424
rect 230 423 231 424
rect 231 423 232 424
rect 232 423 233 424
rect 233 423 234 424
rect 234 423 235 424
rect 235 423 236 424
rect 236 423 237 424
rect 237 423 238 424
rect 238 423 239 424
rect 239 423 240 424
rect 240 423 241 424
rect 241 423 242 424
rect 242 423 243 424
rect 243 423 244 424
rect 244 423 245 424
rect 245 423 246 424
rect 246 423 247 424
rect 247 423 248 424
rect 248 423 249 424
rect 249 423 250 424
rect 250 423 251 424
rect 251 423 252 424
rect 252 423 253 424
rect 253 423 254 424
rect 254 423 255 424
rect 255 423 256 424
rect 256 423 257 424
rect 257 423 258 424
rect 341 423 342 424
rect 342 423 343 424
rect 343 423 344 424
rect 344 423 345 424
rect 345 423 346 424
rect 346 423 347 424
rect 347 423 348 424
rect 348 423 349 424
rect 349 423 350 424
rect 350 423 351 424
rect 351 423 352 424
rect 352 423 353 424
rect 353 423 354 424
rect 360 423 361 424
rect 361 423 362 424
rect 362 423 363 424
rect 363 423 364 424
rect 364 423 365 424
rect 365 423 366 424
rect 366 423 367 424
rect 367 423 368 424
rect 368 423 369 424
rect 369 423 370 424
rect 370 423 371 424
rect 371 423 372 424
rect 372 423 373 424
rect 373 423 374 424
rect 374 423 375 424
rect 375 423 376 424
rect 376 423 377 424
rect 377 423 378 424
rect 158 422 159 423
rect 159 422 160 423
rect 160 422 161 423
rect 221 422 222 423
rect 222 422 223 423
rect 223 422 224 423
rect 224 422 225 423
rect 225 422 226 423
rect 226 422 227 423
rect 227 422 228 423
rect 228 422 229 423
rect 229 422 230 423
rect 230 422 231 423
rect 231 422 232 423
rect 232 422 233 423
rect 233 422 234 423
rect 234 422 235 423
rect 235 422 236 423
rect 236 422 237 423
rect 237 422 238 423
rect 238 422 239 423
rect 239 422 240 423
rect 240 422 241 423
rect 241 422 242 423
rect 242 422 243 423
rect 243 422 244 423
rect 244 422 245 423
rect 245 422 246 423
rect 246 422 247 423
rect 247 422 248 423
rect 248 422 249 423
rect 249 422 250 423
rect 250 422 251 423
rect 251 422 252 423
rect 252 422 253 423
rect 253 422 254 423
rect 254 422 255 423
rect 255 422 256 423
rect 256 422 257 423
rect 257 422 258 423
rect 341 422 342 423
rect 342 422 343 423
rect 343 422 344 423
rect 344 422 345 423
rect 345 422 346 423
rect 346 422 347 423
rect 347 422 348 423
rect 348 422 349 423
rect 349 422 350 423
rect 350 422 351 423
rect 351 422 352 423
rect 352 422 353 423
rect 353 422 354 423
rect 360 422 361 423
rect 361 422 362 423
rect 362 422 363 423
rect 363 422 364 423
rect 364 422 365 423
rect 365 422 366 423
rect 366 422 367 423
rect 367 422 368 423
rect 368 422 369 423
rect 369 422 370 423
rect 370 422 371 423
rect 371 422 372 423
rect 372 422 373 423
rect 373 422 374 423
rect 374 422 375 423
rect 375 422 376 423
rect 154 421 155 422
rect 155 421 156 422
rect 156 421 157 422
rect 157 421 158 422
rect 158 421 159 422
rect 159 421 160 422
rect 160 421 161 422
rect 216 421 217 422
rect 217 421 218 422
rect 218 421 219 422
rect 219 421 220 422
rect 220 421 221 422
rect 221 421 222 422
rect 222 421 223 422
rect 223 421 224 422
rect 224 421 225 422
rect 225 421 226 422
rect 226 421 227 422
rect 227 421 228 422
rect 228 421 229 422
rect 229 421 230 422
rect 230 421 231 422
rect 231 421 232 422
rect 232 421 233 422
rect 233 421 234 422
rect 234 421 235 422
rect 235 421 236 422
rect 236 421 237 422
rect 237 421 238 422
rect 238 421 239 422
rect 239 421 240 422
rect 240 421 241 422
rect 241 421 242 422
rect 242 421 243 422
rect 243 421 244 422
rect 244 421 245 422
rect 245 421 246 422
rect 246 421 247 422
rect 247 421 248 422
rect 248 421 249 422
rect 249 421 250 422
rect 250 421 251 422
rect 251 421 252 422
rect 252 421 253 422
rect 253 421 254 422
rect 254 421 255 422
rect 255 421 256 422
rect 256 421 257 422
rect 257 421 258 422
rect 258 421 259 422
rect 259 421 260 422
rect 260 421 261 422
rect 261 421 262 422
rect 262 421 263 422
rect 263 421 264 422
rect 264 421 265 422
rect 265 421 266 422
rect 266 421 267 422
rect 341 421 342 422
rect 342 421 343 422
rect 343 421 344 422
rect 344 421 345 422
rect 345 421 346 422
rect 346 421 347 422
rect 347 421 348 422
rect 348 421 349 422
rect 349 421 350 422
rect 350 421 351 422
rect 351 421 352 422
rect 352 421 353 422
rect 353 421 354 422
rect 360 421 361 422
rect 361 421 362 422
rect 362 421 363 422
rect 363 421 364 422
rect 364 421 365 422
rect 365 421 366 422
rect 366 421 367 422
rect 367 421 368 422
rect 368 421 369 422
rect 369 421 370 422
rect 370 421 371 422
rect 371 421 372 422
rect 372 421 373 422
rect 373 421 374 422
rect 374 421 375 422
rect 375 421 376 422
rect 154 420 155 421
rect 155 420 156 421
rect 156 420 157 421
rect 157 420 158 421
rect 158 420 159 421
rect 216 420 217 421
rect 217 420 218 421
rect 218 420 219 421
rect 219 420 220 421
rect 220 420 221 421
rect 221 420 222 421
rect 222 420 223 421
rect 223 420 224 421
rect 224 420 225 421
rect 225 420 226 421
rect 226 420 227 421
rect 227 420 228 421
rect 228 420 229 421
rect 229 420 230 421
rect 230 420 231 421
rect 231 420 232 421
rect 232 420 233 421
rect 233 420 234 421
rect 234 420 235 421
rect 235 420 236 421
rect 236 420 237 421
rect 237 420 238 421
rect 238 420 239 421
rect 239 420 240 421
rect 240 420 241 421
rect 241 420 242 421
rect 242 420 243 421
rect 243 420 244 421
rect 244 420 245 421
rect 245 420 246 421
rect 246 420 247 421
rect 247 420 248 421
rect 248 420 249 421
rect 249 420 250 421
rect 250 420 251 421
rect 251 420 252 421
rect 252 420 253 421
rect 253 420 254 421
rect 254 420 255 421
rect 255 420 256 421
rect 256 420 257 421
rect 257 420 258 421
rect 258 420 259 421
rect 259 420 260 421
rect 260 420 261 421
rect 261 420 262 421
rect 262 420 263 421
rect 263 420 264 421
rect 264 420 265 421
rect 265 420 266 421
rect 266 420 267 421
rect 341 420 342 421
rect 342 420 343 421
rect 343 420 344 421
rect 344 420 345 421
rect 345 420 346 421
rect 346 420 347 421
rect 347 420 348 421
rect 348 420 349 421
rect 349 420 350 421
rect 350 420 351 421
rect 351 420 352 421
rect 352 420 353 421
rect 353 420 354 421
rect 360 420 361 421
rect 361 420 362 421
rect 362 420 363 421
rect 363 420 364 421
rect 364 420 365 421
rect 365 420 366 421
rect 366 420 367 421
rect 367 420 368 421
rect 368 420 369 421
rect 369 420 370 421
rect 370 420 371 421
rect 371 420 372 421
rect 372 420 373 421
rect 373 420 374 421
rect 152 419 153 420
rect 153 419 154 420
rect 154 419 155 420
rect 155 419 156 420
rect 156 419 157 420
rect 157 419 158 420
rect 158 419 159 420
rect 210 419 211 420
rect 211 419 212 420
rect 212 419 213 420
rect 213 419 214 420
rect 214 419 215 420
rect 215 419 216 420
rect 216 419 217 420
rect 217 419 218 420
rect 218 419 219 420
rect 219 419 220 420
rect 220 419 221 420
rect 221 419 222 420
rect 222 419 223 420
rect 223 419 224 420
rect 224 419 225 420
rect 225 419 226 420
rect 226 419 227 420
rect 227 419 228 420
rect 228 419 229 420
rect 229 419 230 420
rect 230 419 231 420
rect 231 419 232 420
rect 232 419 233 420
rect 233 419 234 420
rect 234 419 235 420
rect 235 419 236 420
rect 236 419 237 420
rect 237 419 238 420
rect 238 419 239 420
rect 239 419 240 420
rect 240 419 241 420
rect 241 419 242 420
rect 242 419 243 420
rect 243 419 244 420
rect 244 419 245 420
rect 245 419 246 420
rect 246 419 247 420
rect 247 419 248 420
rect 248 419 249 420
rect 249 419 250 420
rect 250 419 251 420
rect 251 419 252 420
rect 252 419 253 420
rect 253 419 254 420
rect 254 419 255 420
rect 255 419 256 420
rect 256 419 257 420
rect 257 419 258 420
rect 258 419 259 420
rect 259 419 260 420
rect 260 419 261 420
rect 261 419 262 420
rect 262 419 263 420
rect 263 419 264 420
rect 264 419 265 420
rect 265 419 266 420
rect 266 419 267 420
rect 267 419 268 420
rect 268 419 269 420
rect 269 419 270 420
rect 270 419 271 420
rect 271 419 272 420
rect 272 419 273 420
rect 273 419 274 420
rect 274 419 275 420
rect 341 419 342 420
rect 342 419 343 420
rect 343 419 344 420
rect 344 419 345 420
rect 345 419 346 420
rect 346 419 347 420
rect 347 419 348 420
rect 348 419 349 420
rect 349 419 350 420
rect 350 419 351 420
rect 351 419 352 420
rect 352 419 353 420
rect 353 419 354 420
rect 360 419 361 420
rect 361 419 362 420
rect 362 419 363 420
rect 363 419 364 420
rect 364 419 365 420
rect 365 419 366 420
rect 366 419 367 420
rect 367 419 368 420
rect 368 419 369 420
rect 369 419 370 420
rect 370 419 371 420
rect 371 419 372 420
rect 372 419 373 420
rect 373 419 374 420
rect 152 418 153 419
rect 153 418 154 419
rect 154 418 155 419
rect 210 418 211 419
rect 211 418 212 419
rect 212 418 213 419
rect 213 418 214 419
rect 214 418 215 419
rect 215 418 216 419
rect 216 418 217 419
rect 217 418 218 419
rect 218 418 219 419
rect 219 418 220 419
rect 220 418 221 419
rect 223 418 224 419
rect 224 418 225 419
rect 225 418 226 419
rect 233 418 234 419
rect 234 418 235 419
rect 235 418 236 419
rect 240 418 241 419
rect 241 418 242 419
rect 242 418 243 419
rect 243 418 244 419
rect 244 418 245 419
rect 246 418 247 419
rect 247 418 248 419
rect 248 418 249 419
rect 249 418 250 419
rect 250 418 251 419
rect 251 418 252 419
rect 252 418 253 419
rect 253 418 254 419
rect 254 418 255 419
rect 255 418 256 419
rect 256 418 257 419
rect 257 418 258 419
rect 258 418 259 419
rect 259 418 260 419
rect 260 418 261 419
rect 261 418 262 419
rect 262 418 263 419
rect 263 418 264 419
rect 264 418 265 419
rect 265 418 266 419
rect 266 418 267 419
rect 267 418 268 419
rect 268 418 269 419
rect 269 418 270 419
rect 270 418 271 419
rect 271 418 272 419
rect 272 418 273 419
rect 273 418 274 419
rect 274 418 275 419
rect 341 418 342 419
rect 342 418 343 419
rect 343 418 344 419
rect 344 418 345 419
rect 345 418 346 419
rect 346 418 347 419
rect 347 418 348 419
rect 348 418 349 419
rect 349 418 350 419
rect 350 418 351 419
rect 351 418 352 419
rect 360 418 361 419
rect 361 418 362 419
rect 362 418 363 419
rect 363 418 364 419
rect 364 418 365 419
rect 365 418 366 419
rect 366 418 367 419
rect 367 418 368 419
rect 368 418 369 419
rect 369 418 370 419
rect 370 418 371 419
rect 371 418 372 419
rect 372 418 373 419
rect 373 418 374 419
rect 150 417 151 418
rect 151 417 152 418
rect 152 417 153 418
rect 153 417 154 418
rect 154 417 155 418
rect 210 417 211 418
rect 211 417 212 418
rect 212 417 213 418
rect 213 417 214 418
rect 214 417 215 418
rect 215 417 216 418
rect 216 417 217 418
rect 217 417 218 418
rect 218 417 219 418
rect 219 417 220 418
rect 220 417 221 418
rect 223 417 224 418
rect 224 417 225 418
rect 225 417 226 418
rect 233 417 234 418
rect 234 417 235 418
rect 235 417 236 418
rect 240 417 241 418
rect 241 417 242 418
rect 242 417 243 418
rect 243 417 244 418
rect 244 417 245 418
rect 246 417 247 418
rect 247 417 248 418
rect 248 417 249 418
rect 249 417 250 418
rect 250 417 251 418
rect 251 417 252 418
rect 252 417 253 418
rect 253 417 254 418
rect 254 417 255 418
rect 255 417 256 418
rect 256 417 257 418
rect 257 417 258 418
rect 258 417 259 418
rect 259 417 260 418
rect 260 417 261 418
rect 261 417 262 418
rect 262 417 263 418
rect 263 417 264 418
rect 264 417 265 418
rect 265 417 266 418
rect 266 417 267 418
rect 267 417 268 418
rect 268 417 269 418
rect 269 417 270 418
rect 270 417 271 418
rect 271 417 272 418
rect 272 417 273 418
rect 273 417 274 418
rect 274 417 275 418
rect 275 417 276 418
rect 276 417 277 418
rect 277 417 278 418
rect 278 417 279 418
rect 279 417 280 418
rect 280 417 281 418
rect 281 417 282 418
rect 339 417 340 418
rect 340 417 341 418
rect 341 417 342 418
rect 342 417 343 418
rect 343 417 344 418
rect 344 417 345 418
rect 345 417 346 418
rect 346 417 347 418
rect 347 417 348 418
rect 348 417 349 418
rect 349 417 350 418
rect 350 417 351 418
rect 351 417 352 418
rect 352 417 353 418
rect 353 417 354 418
rect 358 417 359 418
rect 359 417 360 418
rect 360 417 361 418
rect 361 417 362 418
rect 362 417 363 418
rect 363 417 364 418
rect 364 417 365 418
rect 365 417 366 418
rect 366 417 367 418
rect 367 417 368 418
rect 368 417 369 418
rect 369 417 370 418
rect 370 417 371 418
rect 371 417 372 418
rect 372 417 373 418
rect 373 417 374 418
rect 150 416 151 417
rect 151 416 152 417
rect 152 416 153 417
rect 257 416 258 417
rect 258 416 259 417
rect 259 416 260 417
rect 260 416 261 417
rect 261 416 262 417
rect 262 416 263 417
rect 263 416 264 417
rect 264 416 265 417
rect 265 416 266 417
rect 266 416 267 417
rect 267 416 268 417
rect 268 416 269 417
rect 269 416 270 417
rect 270 416 271 417
rect 271 416 272 417
rect 272 416 273 417
rect 273 416 274 417
rect 274 416 275 417
rect 275 416 276 417
rect 276 416 277 417
rect 277 416 278 417
rect 278 416 279 417
rect 279 416 280 417
rect 280 416 281 417
rect 281 416 282 417
rect 339 416 340 417
rect 340 416 341 417
rect 341 416 342 417
rect 342 416 343 417
rect 343 416 344 417
rect 344 416 345 417
rect 345 416 346 417
rect 346 416 347 417
rect 347 416 348 417
rect 348 416 349 417
rect 349 416 350 417
rect 350 416 351 417
rect 351 416 352 417
rect 352 416 353 417
rect 353 416 354 417
rect 358 416 359 417
rect 359 416 360 417
rect 360 416 361 417
rect 361 416 362 417
rect 362 416 363 417
rect 363 416 364 417
rect 364 416 365 417
rect 365 416 366 417
rect 366 416 367 417
rect 367 416 368 417
rect 368 416 369 417
rect 369 416 370 417
rect 370 416 371 417
rect 371 416 372 417
rect 147 415 148 416
rect 148 415 149 416
rect 149 415 150 416
rect 150 415 151 416
rect 151 415 152 416
rect 152 415 153 416
rect 257 415 258 416
rect 258 415 259 416
rect 259 415 260 416
rect 260 415 261 416
rect 261 415 262 416
rect 262 415 263 416
rect 263 415 264 416
rect 264 415 265 416
rect 265 415 266 416
rect 266 415 267 416
rect 267 415 268 416
rect 268 415 269 416
rect 269 415 270 416
rect 270 415 271 416
rect 271 415 272 416
rect 272 415 273 416
rect 273 415 274 416
rect 274 415 275 416
rect 275 415 276 416
rect 276 415 277 416
rect 277 415 278 416
rect 278 415 279 416
rect 279 415 280 416
rect 280 415 281 416
rect 281 415 282 416
rect 282 415 283 416
rect 283 415 284 416
rect 284 415 285 416
rect 285 415 286 416
rect 339 415 340 416
rect 340 415 341 416
rect 341 415 342 416
rect 342 415 343 416
rect 343 415 344 416
rect 344 415 345 416
rect 345 415 346 416
rect 346 415 347 416
rect 347 415 348 416
rect 348 415 349 416
rect 349 415 350 416
rect 350 415 351 416
rect 351 415 352 416
rect 352 415 353 416
rect 353 415 354 416
rect 356 415 357 416
rect 357 415 358 416
rect 358 415 359 416
rect 359 415 360 416
rect 360 415 361 416
rect 361 415 362 416
rect 362 415 363 416
rect 363 415 364 416
rect 364 415 365 416
rect 365 415 366 416
rect 366 415 367 416
rect 367 415 368 416
rect 368 415 369 416
rect 369 415 370 416
rect 370 415 371 416
rect 371 415 372 416
rect 147 414 148 415
rect 148 414 149 415
rect 149 414 150 415
rect 150 414 151 415
rect 266 414 267 415
rect 267 414 268 415
rect 268 414 269 415
rect 269 414 270 415
rect 270 414 271 415
rect 271 414 272 415
rect 272 414 273 415
rect 273 414 274 415
rect 274 414 275 415
rect 275 414 276 415
rect 276 414 277 415
rect 277 414 278 415
rect 278 414 279 415
rect 279 414 280 415
rect 280 414 281 415
rect 281 414 282 415
rect 282 414 283 415
rect 283 414 284 415
rect 284 414 285 415
rect 285 414 286 415
rect 341 414 342 415
rect 342 414 343 415
rect 343 414 344 415
rect 344 414 345 415
rect 345 414 346 415
rect 346 414 347 415
rect 347 414 348 415
rect 348 414 349 415
rect 349 414 350 415
rect 350 414 351 415
rect 351 414 352 415
rect 356 414 357 415
rect 357 414 358 415
rect 358 414 359 415
rect 359 414 360 415
rect 360 414 361 415
rect 361 414 362 415
rect 362 414 363 415
rect 363 414 364 415
rect 364 414 365 415
rect 365 414 366 415
rect 366 414 367 415
rect 367 414 368 415
rect 368 414 369 415
rect 369 414 370 415
rect 143 413 144 414
rect 144 413 145 414
rect 145 413 146 414
rect 146 413 147 414
rect 147 413 148 414
rect 148 413 149 414
rect 149 413 150 414
rect 150 413 151 414
rect 199 413 200 414
rect 200 413 201 414
rect 201 413 202 414
rect 266 413 267 414
rect 267 413 268 414
rect 268 413 269 414
rect 269 413 270 414
rect 270 413 271 414
rect 271 413 272 414
rect 272 413 273 414
rect 273 413 274 414
rect 274 413 275 414
rect 275 413 276 414
rect 276 413 277 414
rect 277 413 278 414
rect 278 413 279 414
rect 279 413 280 414
rect 280 413 281 414
rect 281 413 282 414
rect 282 413 283 414
rect 283 413 284 414
rect 284 413 285 414
rect 285 413 286 414
rect 286 413 287 414
rect 287 413 288 414
rect 288 413 289 414
rect 289 413 290 414
rect 290 413 291 414
rect 291 413 292 414
rect 341 413 342 414
rect 342 413 343 414
rect 343 413 344 414
rect 344 413 345 414
rect 345 413 346 414
rect 346 413 347 414
rect 347 413 348 414
rect 348 413 349 414
rect 349 413 350 414
rect 350 413 351 414
rect 351 413 352 414
rect 356 413 357 414
rect 357 413 358 414
rect 358 413 359 414
rect 359 413 360 414
rect 360 413 361 414
rect 361 413 362 414
rect 362 413 363 414
rect 363 413 364 414
rect 364 413 365 414
rect 365 413 366 414
rect 366 413 367 414
rect 367 413 368 414
rect 368 413 369 414
rect 369 413 370 414
rect 143 412 144 413
rect 144 412 145 413
rect 145 412 146 413
rect 146 412 147 413
rect 147 412 148 413
rect 148 412 149 413
rect 199 412 200 413
rect 200 412 201 413
rect 201 412 202 413
rect 274 412 275 413
rect 275 412 276 413
rect 276 412 277 413
rect 277 412 278 413
rect 278 412 279 413
rect 279 412 280 413
rect 280 412 281 413
rect 281 412 282 413
rect 282 412 283 413
rect 283 412 284 413
rect 284 412 285 413
rect 285 412 286 413
rect 286 412 287 413
rect 287 412 288 413
rect 288 412 289 413
rect 289 412 290 413
rect 290 412 291 413
rect 291 412 292 413
rect 341 412 342 413
rect 342 412 343 413
rect 343 412 344 413
rect 344 412 345 413
rect 345 412 346 413
rect 346 412 347 413
rect 347 412 348 413
rect 348 412 349 413
rect 349 412 350 413
rect 350 412 351 413
rect 351 412 352 413
rect 356 412 357 413
rect 357 412 358 413
rect 358 412 359 413
rect 359 412 360 413
rect 360 412 361 413
rect 361 412 362 413
rect 362 412 363 413
rect 363 412 364 413
rect 364 412 365 413
rect 365 412 366 413
rect 366 412 367 413
rect 367 412 368 413
rect 368 412 369 413
rect 369 412 370 413
rect 141 411 142 412
rect 142 411 143 412
rect 143 411 144 412
rect 144 411 145 412
rect 145 411 146 412
rect 146 411 147 412
rect 147 411 148 412
rect 148 411 149 412
rect 195 411 196 412
rect 196 411 197 412
rect 197 411 198 412
rect 198 411 199 412
rect 199 411 200 412
rect 200 411 201 412
rect 201 411 202 412
rect 274 411 275 412
rect 275 411 276 412
rect 276 411 277 412
rect 277 411 278 412
rect 278 411 279 412
rect 279 411 280 412
rect 280 411 281 412
rect 281 411 282 412
rect 282 411 283 412
rect 283 411 284 412
rect 284 411 285 412
rect 285 411 286 412
rect 286 411 287 412
rect 287 411 288 412
rect 288 411 289 412
rect 289 411 290 412
rect 290 411 291 412
rect 291 411 292 412
rect 292 411 293 412
rect 293 411 294 412
rect 294 411 295 412
rect 295 411 296 412
rect 296 411 297 412
rect 339 411 340 412
rect 340 411 341 412
rect 341 411 342 412
rect 342 411 343 412
rect 343 411 344 412
rect 344 411 345 412
rect 345 411 346 412
rect 346 411 347 412
rect 347 411 348 412
rect 348 411 349 412
rect 349 411 350 412
rect 350 411 351 412
rect 351 411 352 412
rect 356 411 357 412
rect 357 411 358 412
rect 358 411 359 412
rect 359 411 360 412
rect 360 411 361 412
rect 361 411 362 412
rect 362 411 363 412
rect 363 411 364 412
rect 364 411 365 412
rect 365 411 366 412
rect 366 411 367 412
rect 367 411 368 412
rect 368 411 369 412
rect 369 411 370 412
rect 141 410 142 411
rect 142 410 143 411
rect 143 410 144 411
rect 144 410 145 411
rect 145 410 146 411
rect 195 410 196 411
rect 196 410 197 411
rect 197 410 198 411
rect 198 410 199 411
rect 199 410 200 411
rect 281 410 282 411
rect 282 410 283 411
rect 283 410 284 411
rect 284 410 285 411
rect 285 410 286 411
rect 286 410 287 411
rect 287 410 288 411
rect 288 410 289 411
rect 289 410 290 411
rect 290 410 291 411
rect 291 410 292 411
rect 292 410 293 411
rect 293 410 294 411
rect 294 410 295 411
rect 295 410 296 411
rect 296 410 297 411
rect 339 410 340 411
rect 340 410 341 411
rect 341 410 342 411
rect 342 410 343 411
rect 343 410 344 411
rect 344 410 345 411
rect 345 410 346 411
rect 346 410 347 411
rect 347 410 348 411
rect 348 410 349 411
rect 349 410 350 411
rect 350 410 351 411
rect 351 410 352 411
rect 356 410 357 411
rect 357 410 358 411
rect 358 410 359 411
rect 359 410 360 411
rect 360 410 361 411
rect 361 410 362 411
rect 362 410 363 411
rect 363 410 364 411
rect 364 410 365 411
rect 365 410 366 411
rect 366 410 367 411
rect 367 410 368 411
rect 368 410 369 411
rect 137 409 138 410
rect 138 409 139 410
rect 139 409 140 410
rect 140 409 141 410
rect 141 409 142 410
rect 142 409 143 410
rect 143 409 144 410
rect 144 409 145 410
rect 145 409 146 410
rect 191 409 192 410
rect 192 409 193 410
rect 193 409 194 410
rect 194 409 195 410
rect 195 409 196 410
rect 196 409 197 410
rect 197 409 198 410
rect 198 409 199 410
rect 199 409 200 410
rect 281 409 282 410
rect 282 409 283 410
rect 283 409 284 410
rect 284 409 285 410
rect 285 409 286 410
rect 286 409 287 410
rect 287 409 288 410
rect 288 409 289 410
rect 289 409 290 410
rect 290 409 291 410
rect 291 409 292 410
rect 292 409 293 410
rect 293 409 294 410
rect 294 409 295 410
rect 295 409 296 410
rect 296 409 297 410
rect 297 409 298 410
rect 298 409 299 410
rect 299 409 300 410
rect 300 409 301 410
rect 301 409 302 410
rect 302 409 303 410
rect 339 409 340 410
rect 340 409 341 410
rect 341 409 342 410
rect 342 409 343 410
rect 343 409 344 410
rect 344 409 345 410
rect 345 409 346 410
rect 346 409 347 410
rect 347 409 348 410
rect 348 409 349 410
rect 349 409 350 410
rect 350 409 351 410
rect 351 409 352 410
rect 354 409 355 410
rect 355 409 356 410
rect 356 409 357 410
rect 357 409 358 410
rect 358 409 359 410
rect 359 409 360 410
rect 360 409 361 410
rect 361 409 362 410
rect 362 409 363 410
rect 363 409 364 410
rect 364 409 365 410
rect 365 409 366 410
rect 366 409 367 410
rect 367 409 368 410
rect 368 409 369 410
rect 137 408 138 409
rect 138 408 139 409
rect 139 408 140 409
rect 140 408 141 409
rect 141 408 142 409
rect 142 408 143 409
rect 143 408 144 409
rect 191 408 192 409
rect 192 408 193 409
rect 193 408 194 409
rect 194 408 195 409
rect 195 408 196 409
rect 196 408 197 409
rect 197 408 198 409
rect 289 408 290 409
rect 290 408 291 409
rect 291 408 292 409
rect 292 408 293 409
rect 293 408 294 409
rect 294 408 295 409
rect 295 408 296 409
rect 296 408 297 409
rect 297 408 298 409
rect 298 408 299 409
rect 299 408 300 409
rect 300 408 301 409
rect 301 408 302 409
rect 302 408 303 409
rect 341 408 342 409
rect 342 408 343 409
rect 343 408 344 409
rect 344 408 345 409
rect 345 408 346 409
rect 346 408 347 409
rect 347 408 348 409
rect 348 408 349 409
rect 349 408 350 409
rect 350 408 351 409
rect 351 408 352 409
rect 354 408 355 409
rect 355 408 356 409
rect 356 408 357 409
rect 357 408 358 409
rect 358 408 359 409
rect 359 408 360 409
rect 360 408 361 409
rect 361 408 362 409
rect 362 408 363 409
rect 363 408 364 409
rect 364 408 365 409
rect 365 408 366 409
rect 366 408 367 409
rect 367 408 368 409
rect 368 408 369 409
rect 135 407 136 408
rect 136 407 137 408
rect 137 407 138 408
rect 138 407 139 408
rect 139 407 140 408
rect 140 407 141 408
rect 141 407 142 408
rect 142 407 143 408
rect 143 407 144 408
rect 188 407 189 408
rect 189 407 190 408
rect 190 407 191 408
rect 191 407 192 408
rect 192 407 193 408
rect 193 407 194 408
rect 194 407 195 408
rect 195 407 196 408
rect 196 407 197 408
rect 197 407 198 408
rect 289 407 290 408
rect 290 407 291 408
rect 291 407 292 408
rect 292 407 293 408
rect 293 407 294 408
rect 294 407 295 408
rect 295 407 296 408
rect 296 407 297 408
rect 297 407 298 408
rect 298 407 299 408
rect 299 407 300 408
rect 300 407 301 408
rect 301 407 302 408
rect 302 407 303 408
rect 303 407 304 408
rect 304 407 305 408
rect 305 407 306 408
rect 306 407 307 408
rect 341 407 342 408
rect 342 407 343 408
rect 343 407 344 408
rect 344 407 345 408
rect 345 407 346 408
rect 346 407 347 408
rect 347 407 348 408
rect 348 407 349 408
rect 349 407 350 408
rect 350 407 351 408
rect 351 407 352 408
rect 354 407 355 408
rect 355 407 356 408
rect 356 407 357 408
rect 357 407 358 408
rect 358 407 359 408
rect 359 407 360 408
rect 360 407 361 408
rect 361 407 362 408
rect 362 407 363 408
rect 363 407 364 408
rect 364 407 365 408
rect 365 407 366 408
rect 366 407 367 408
rect 367 407 368 408
rect 368 407 369 408
rect 135 406 136 407
rect 136 406 137 407
rect 137 406 138 407
rect 138 406 139 407
rect 139 406 140 407
rect 140 406 141 407
rect 141 406 142 407
rect 188 406 189 407
rect 189 406 190 407
rect 190 406 191 407
rect 191 406 192 407
rect 192 406 193 407
rect 193 406 194 407
rect 194 406 195 407
rect 195 406 196 407
rect 196 406 197 407
rect 197 406 198 407
rect 296 406 297 407
rect 297 406 298 407
rect 298 406 299 407
rect 299 406 300 407
rect 300 406 301 407
rect 301 406 302 407
rect 302 406 303 407
rect 303 406 304 407
rect 304 406 305 407
rect 305 406 306 407
rect 306 406 307 407
rect 341 406 342 407
rect 342 406 343 407
rect 343 406 344 407
rect 344 406 345 407
rect 345 406 346 407
rect 346 406 347 407
rect 347 406 348 407
rect 348 406 349 407
rect 349 406 350 407
rect 350 406 351 407
rect 351 406 352 407
rect 356 406 357 407
rect 357 406 358 407
rect 358 406 359 407
rect 359 406 360 407
rect 360 406 361 407
rect 361 406 362 407
rect 362 406 363 407
rect 363 406 364 407
rect 364 406 365 407
rect 365 406 366 407
rect 366 406 367 407
rect 132 405 133 406
rect 133 405 134 406
rect 134 405 135 406
rect 135 405 136 406
rect 136 405 137 406
rect 137 405 138 406
rect 138 405 139 406
rect 139 405 140 406
rect 140 405 141 406
rect 141 405 142 406
rect 186 405 187 406
rect 187 405 188 406
rect 188 405 189 406
rect 189 405 190 406
rect 190 405 191 406
rect 191 405 192 406
rect 192 405 193 406
rect 193 405 194 406
rect 194 405 195 406
rect 195 405 196 406
rect 196 405 197 406
rect 197 405 198 406
rect 296 405 297 406
rect 297 405 298 406
rect 298 405 299 406
rect 299 405 300 406
rect 300 405 301 406
rect 301 405 302 406
rect 302 405 303 406
rect 303 405 304 406
rect 304 405 305 406
rect 305 405 306 406
rect 306 405 307 406
rect 307 405 308 406
rect 308 405 309 406
rect 309 405 310 406
rect 310 405 311 406
rect 311 405 312 406
rect 341 405 342 406
rect 342 405 343 406
rect 343 405 344 406
rect 344 405 345 406
rect 345 405 346 406
rect 346 405 347 406
rect 347 405 348 406
rect 348 405 349 406
rect 349 405 350 406
rect 350 405 351 406
rect 351 405 352 406
rect 354 405 355 406
rect 355 405 356 406
rect 356 405 357 406
rect 357 405 358 406
rect 358 405 359 406
rect 359 405 360 406
rect 360 405 361 406
rect 361 405 362 406
rect 362 405 363 406
rect 363 405 364 406
rect 364 405 365 406
rect 365 405 366 406
rect 366 405 367 406
rect 367 405 368 406
rect 368 405 369 406
rect 132 404 133 405
rect 133 404 134 405
rect 134 404 135 405
rect 135 404 136 405
rect 136 404 137 405
rect 137 404 138 405
rect 186 404 187 405
rect 187 404 188 405
rect 188 404 189 405
rect 189 404 190 405
rect 190 404 191 405
rect 191 404 192 405
rect 192 404 193 405
rect 193 404 194 405
rect 194 404 195 405
rect 195 404 196 405
rect 302 404 303 405
rect 303 404 304 405
rect 304 404 305 405
rect 305 404 306 405
rect 306 404 307 405
rect 307 404 308 405
rect 308 404 309 405
rect 309 404 310 405
rect 310 404 311 405
rect 311 404 312 405
rect 341 404 342 405
rect 342 404 343 405
rect 343 404 344 405
rect 344 404 345 405
rect 345 404 346 405
rect 346 404 347 405
rect 347 404 348 405
rect 348 404 349 405
rect 349 404 350 405
rect 350 404 351 405
rect 351 404 352 405
rect 354 404 355 405
rect 355 404 356 405
rect 356 404 357 405
rect 357 404 358 405
rect 358 404 359 405
rect 359 404 360 405
rect 360 404 361 405
rect 361 404 362 405
rect 362 404 363 405
rect 363 404 364 405
rect 364 404 365 405
rect 365 404 366 405
rect 366 404 367 405
rect 367 404 368 405
rect 368 404 369 405
rect 128 403 129 404
rect 129 403 130 404
rect 130 403 131 404
rect 131 403 132 404
rect 132 403 133 404
rect 133 403 134 404
rect 134 403 135 404
rect 135 403 136 404
rect 136 403 137 404
rect 137 403 138 404
rect 182 403 183 404
rect 183 403 184 404
rect 184 403 185 404
rect 185 403 186 404
rect 186 403 187 404
rect 187 403 188 404
rect 188 403 189 404
rect 189 403 190 404
rect 190 403 191 404
rect 191 403 192 404
rect 192 403 193 404
rect 193 403 194 404
rect 194 403 195 404
rect 195 403 196 404
rect 302 403 303 404
rect 303 403 304 404
rect 304 403 305 404
rect 305 403 306 404
rect 306 403 307 404
rect 307 403 308 404
rect 308 403 309 404
rect 309 403 310 404
rect 310 403 311 404
rect 311 403 312 404
rect 312 403 313 404
rect 313 403 314 404
rect 314 403 315 404
rect 315 403 316 404
rect 316 403 317 404
rect 317 403 318 404
rect 339 403 340 404
rect 340 403 341 404
rect 341 403 342 404
rect 342 403 343 404
rect 343 403 344 404
rect 344 403 345 404
rect 345 403 346 404
rect 346 403 347 404
rect 347 403 348 404
rect 348 403 349 404
rect 349 403 350 404
rect 350 403 351 404
rect 351 403 352 404
rect 354 403 355 404
rect 355 403 356 404
rect 356 403 357 404
rect 357 403 358 404
rect 358 403 359 404
rect 359 403 360 404
rect 360 403 361 404
rect 361 403 362 404
rect 362 403 363 404
rect 363 403 364 404
rect 364 403 365 404
rect 365 403 366 404
rect 366 403 367 404
rect 367 403 368 404
rect 368 403 369 404
rect 128 402 129 403
rect 129 402 130 403
rect 130 402 131 403
rect 131 402 132 403
rect 132 402 133 403
rect 133 402 134 403
rect 134 402 135 403
rect 135 402 136 403
rect 182 402 183 403
rect 183 402 184 403
rect 184 402 185 403
rect 185 402 186 403
rect 186 402 187 403
rect 187 402 188 403
rect 188 402 189 403
rect 189 402 190 403
rect 190 402 191 403
rect 191 402 192 403
rect 192 402 193 403
rect 193 402 194 403
rect 309 402 310 403
rect 310 402 311 403
rect 311 402 312 403
rect 312 402 313 403
rect 313 402 314 403
rect 314 402 315 403
rect 315 402 316 403
rect 316 402 317 403
rect 317 402 318 403
rect 339 402 340 403
rect 340 402 341 403
rect 341 402 342 403
rect 342 402 343 403
rect 343 402 344 403
rect 344 402 345 403
rect 345 402 346 403
rect 346 402 347 403
rect 347 402 348 403
rect 348 402 349 403
rect 349 402 350 403
rect 354 402 355 403
rect 355 402 356 403
rect 356 402 357 403
rect 357 402 358 403
rect 358 402 359 403
rect 359 402 360 403
rect 360 402 361 403
rect 361 402 362 403
rect 362 402 363 403
rect 363 402 364 403
rect 364 402 365 403
rect 365 402 366 403
rect 366 402 367 403
rect 124 401 125 402
rect 125 401 126 402
rect 126 401 127 402
rect 127 401 128 402
rect 128 401 129 402
rect 129 401 130 402
rect 130 401 131 402
rect 131 401 132 402
rect 132 401 133 402
rect 133 401 134 402
rect 134 401 135 402
rect 135 401 136 402
rect 180 401 181 402
rect 181 401 182 402
rect 182 401 183 402
rect 183 401 184 402
rect 184 401 185 402
rect 185 401 186 402
rect 186 401 187 402
rect 187 401 188 402
rect 188 401 189 402
rect 189 401 190 402
rect 190 401 191 402
rect 191 401 192 402
rect 192 401 193 402
rect 193 401 194 402
rect 309 401 310 402
rect 310 401 311 402
rect 311 401 312 402
rect 312 401 313 402
rect 313 401 314 402
rect 314 401 315 402
rect 315 401 316 402
rect 316 401 317 402
rect 317 401 318 402
rect 318 401 319 402
rect 319 401 320 402
rect 320 401 321 402
rect 321 401 322 402
rect 339 401 340 402
rect 340 401 341 402
rect 341 401 342 402
rect 342 401 343 402
rect 343 401 344 402
rect 344 401 345 402
rect 345 401 346 402
rect 346 401 347 402
rect 347 401 348 402
rect 348 401 349 402
rect 349 401 350 402
rect 350 401 351 402
rect 351 401 352 402
rect 354 401 355 402
rect 355 401 356 402
rect 356 401 357 402
rect 357 401 358 402
rect 358 401 359 402
rect 359 401 360 402
rect 360 401 361 402
rect 361 401 362 402
rect 362 401 363 402
rect 363 401 364 402
rect 364 401 365 402
rect 365 401 366 402
rect 366 401 367 402
rect 367 401 368 402
rect 368 401 369 402
rect 124 400 125 401
rect 125 400 126 401
rect 126 400 127 401
rect 127 400 128 401
rect 128 400 129 401
rect 129 400 130 401
rect 130 400 131 401
rect 131 400 132 401
rect 132 400 133 401
rect 180 400 181 401
rect 181 400 182 401
rect 182 400 183 401
rect 183 400 184 401
rect 184 400 185 401
rect 185 400 186 401
rect 186 400 187 401
rect 187 400 188 401
rect 188 400 189 401
rect 189 400 190 401
rect 190 400 191 401
rect 191 400 192 401
rect 315 400 316 401
rect 316 400 317 401
rect 317 400 318 401
rect 318 400 319 401
rect 319 400 320 401
rect 320 400 321 401
rect 321 400 322 401
rect 341 400 342 401
rect 342 400 343 401
rect 343 400 344 401
rect 344 400 345 401
rect 345 400 346 401
rect 346 400 347 401
rect 347 400 348 401
rect 348 400 349 401
rect 349 400 350 401
rect 350 400 351 401
rect 351 400 352 401
rect 354 400 355 401
rect 355 400 356 401
rect 356 400 357 401
rect 357 400 358 401
rect 358 400 359 401
rect 359 400 360 401
rect 360 400 361 401
rect 361 400 362 401
rect 362 400 363 401
rect 363 400 364 401
rect 364 400 365 401
rect 365 400 366 401
rect 366 400 367 401
rect 367 400 368 401
rect 368 400 369 401
rect 122 399 123 400
rect 123 399 124 400
rect 124 399 125 400
rect 125 399 126 400
rect 126 399 127 400
rect 127 399 128 400
rect 128 399 129 400
rect 129 399 130 400
rect 130 399 131 400
rect 131 399 132 400
rect 132 399 133 400
rect 176 399 177 400
rect 177 399 178 400
rect 178 399 179 400
rect 179 399 180 400
rect 180 399 181 400
rect 181 399 182 400
rect 182 399 183 400
rect 183 399 184 400
rect 184 399 185 400
rect 185 399 186 400
rect 186 399 187 400
rect 187 399 188 400
rect 188 399 189 400
rect 189 399 190 400
rect 190 399 191 400
rect 191 399 192 400
rect 315 399 316 400
rect 316 399 317 400
rect 317 399 318 400
rect 318 399 319 400
rect 319 399 320 400
rect 320 399 321 400
rect 321 399 322 400
rect 323 399 324 400
rect 324 399 325 400
rect 339 399 340 400
rect 340 399 341 400
rect 341 399 342 400
rect 342 399 343 400
rect 343 399 344 400
rect 344 399 345 400
rect 345 399 346 400
rect 346 399 347 400
rect 347 399 348 400
rect 348 399 349 400
rect 349 399 350 400
rect 350 399 351 400
rect 351 399 352 400
rect 354 399 355 400
rect 355 399 356 400
rect 356 399 357 400
rect 357 399 358 400
rect 358 399 359 400
rect 359 399 360 400
rect 360 399 361 400
rect 361 399 362 400
rect 362 399 363 400
rect 363 399 364 400
rect 364 399 365 400
rect 365 399 366 400
rect 366 399 367 400
rect 367 399 368 400
rect 368 399 369 400
rect 394 399 395 400
rect 395 399 396 400
rect 396 399 397 400
rect 444 399 445 400
rect 445 399 446 400
rect 446 399 447 400
rect 452 399 453 400
rect 453 399 454 400
rect 454 399 455 400
rect 457 399 458 400
rect 458 399 459 400
rect 459 399 460 400
rect 122 398 123 399
rect 123 398 124 399
rect 124 398 125 399
rect 125 398 126 399
rect 126 398 127 399
rect 127 398 128 399
rect 128 398 129 399
rect 129 398 130 399
rect 130 398 131 399
rect 176 398 177 399
rect 177 398 178 399
rect 178 398 179 399
rect 179 398 180 399
rect 180 398 181 399
rect 181 398 182 399
rect 182 398 183 399
rect 183 398 184 399
rect 184 398 185 399
rect 185 398 186 399
rect 186 398 187 399
rect 187 398 188 399
rect 188 398 189 399
rect 189 398 190 399
rect 190 398 191 399
rect 323 398 324 399
rect 324 398 325 399
rect 339 398 340 399
rect 340 398 341 399
rect 341 398 342 399
rect 342 398 343 399
rect 343 398 344 399
rect 344 398 345 399
rect 345 398 346 399
rect 346 398 347 399
rect 347 398 348 399
rect 348 398 349 399
rect 349 398 350 399
rect 350 398 351 399
rect 351 398 352 399
rect 354 398 355 399
rect 355 398 356 399
rect 356 398 357 399
rect 357 398 358 399
rect 358 398 359 399
rect 359 398 360 399
rect 360 398 361 399
rect 361 398 362 399
rect 362 398 363 399
rect 363 398 364 399
rect 364 398 365 399
rect 365 398 366 399
rect 366 398 367 399
rect 367 398 368 399
rect 368 398 369 399
rect 394 398 395 399
rect 395 398 396 399
rect 396 398 397 399
rect 444 398 445 399
rect 445 398 446 399
rect 446 398 447 399
rect 452 398 453 399
rect 453 398 454 399
rect 454 398 455 399
rect 457 398 458 399
rect 458 398 459 399
rect 459 398 460 399
rect 118 397 119 398
rect 119 397 120 398
rect 120 397 121 398
rect 121 397 122 398
rect 122 397 123 398
rect 123 397 124 398
rect 124 397 125 398
rect 125 397 126 398
rect 126 397 127 398
rect 127 397 128 398
rect 128 397 129 398
rect 129 397 130 398
rect 130 397 131 398
rect 175 397 176 398
rect 176 397 177 398
rect 177 397 178 398
rect 178 397 179 398
rect 179 397 180 398
rect 180 397 181 398
rect 181 397 182 398
rect 182 397 183 398
rect 183 397 184 398
rect 184 397 185 398
rect 185 397 186 398
rect 186 397 187 398
rect 187 397 188 398
rect 188 397 189 398
rect 189 397 190 398
rect 190 397 191 398
rect 323 397 324 398
rect 324 397 325 398
rect 339 397 340 398
rect 340 397 341 398
rect 341 397 342 398
rect 342 397 343 398
rect 343 397 344 398
rect 344 397 345 398
rect 345 397 346 398
rect 346 397 347 398
rect 347 397 348 398
rect 348 397 349 398
rect 349 397 350 398
rect 350 397 351 398
rect 351 397 352 398
rect 354 397 355 398
rect 355 397 356 398
rect 356 397 357 398
rect 357 397 358 398
rect 358 397 359 398
rect 359 397 360 398
rect 360 397 361 398
rect 361 397 362 398
rect 362 397 363 398
rect 363 397 364 398
rect 364 397 365 398
rect 365 397 366 398
rect 366 397 367 398
rect 367 397 368 398
rect 368 397 369 398
rect 386 397 387 398
rect 387 397 388 398
rect 388 397 389 398
rect 389 397 390 398
rect 390 397 391 398
rect 391 397 392 398
rect 392 397 393 398
rect 393 397 394 398
rect 394 397 395 398
rect 395 397 396 398
rect 396 397 397 398
rect 397 397 398 398
rect 398 397 399 398
rect 399 397 400 398
rect 400 397 401 398
rect 401 397 402 398
rect 402 397 403 398
rect 403 397 404 398
rect 404 397 405 398
rect 405 397 406 398
rect 406 397 407 398
rect 407 397 408 398
rect 408 397 409 398
rect 409 397 410 398
rect 410 397 411 398
rect 411 397 412 398
rect 412 397 413 398
rect 413 397 414 398
rect 414 397 415 398
rect 415 397 416 398
rect 416 397 417 398
rect 417 397 418 398
rect 418 397 419 398
rect 419 397 420 398
rect 420 397 421 398
rect 421 397 422 398
rect 422 397 423 398
rect 423 397 424 398
rect 424 397 425 398
rect 425 397 426 398
rect 426 397 427 398
rect 427 397 428 398
rect 428 397 429 398
rect 429 397 430 398
rect 430 397 431 398
rect 431 397 432 398
rect 432 397 433 398
rect 433 397 434 398
rect 434 397 435 398
rect 435 397 436 398
rect 436 397 437 398
rect 437 397 438 398
rect 438 397 439 398
rect 439 397 440 398
rect 440 397 441 398
rect 441 397 442 398
rect 442 397 443 398
rect 443 397 444 398
rect 444 397 445 398
rect 445 397 446 398
rect 446 397 447 398
rect 447 397 448 398
rect 448 397 449 398
rect 449 397 450 398
rect 450 397 451 398
rect 451 397 452 398
rect 452 397 453 398
rect 453 397 454 398
rect 454 397 455 398
rect 455 397 456 398
rect 456 397 457 398
rect 457 397 458 398
rect 458 397 459 398
rect 459 397 460 398
rect 460 397 461 398
rect 461 397 462 398
rect 462 397 463 398
rect 463 397 464 398
rect 464 397 465 398
rect 465 397 466 398
rect 466 397 467 398
rect 467 397 468 398
rect 468 397 469 398
rect 469 397 470 398
rect 470 397 471 398
rect 471 397 472 398
rect 472 397 473 398
rect 473 397 474 398
rect 474 397 475 398
rect 476 397 477 398
rect 477 397 478 398
rect 478 397 479 398
rect 118 396 119 397
rect 119 396 120 397
rect 120 396 121 397
rect 121 396 122 397
rect 122 396 123 397
rect 123 396 124 397
rect 124 396 125 397
rect 125 396 126 397
rect 126 396 127 397
rect 127 396 128 397
rect 128 396 129 397
rect 175 396 176 397
rect 176 396 177 397
rect 177 396 178 397
rect 178 396 179 397
rect 179 396 180 397
rect 180 396 181 397
rect 181 396 182 397
rect 182 396 183 397
rect 183 396 184 397
rect 184 396 185 397
rect 185 396 186 397
rect 186 396 187 397
rect 187 396 188 397
rect 188 396 189 397
rect 341 396 342 397
rect 342 396 343 397
rect 343 396 344 397
rect 344 396 345 397
rect 345 396 346 397
rect 346 396 347 397
rect 347 396 348 397
rect 348 396 349 397
rect 349 396 350 397
rect 354 396 355 397
rect 355 396 356 397
rect 356 396 357 397
rect 357 396 358 397
rect 358 396 359 397
rect 359 396 360 397
rect 360 396 361 397
rect 361 396 362 397
rect 362 396 363 397
rect 363 396 364 397
rect 364 396 365 397
rect 365 396 366 397
rect 366 396 367 397
rect 386 396 387 397
rect 387 396 388 397
rect 388 396 389 397
rect 389 396 390 397
rect 390 396 391 397
rect 391 396 392 397
rect 392 396 393 397
rect 393 396 394 397
rect 394 396 395 397
rect 395 396 396 397
rect 396 396 397 397
rect 397 396 398 397
rect 398 396 399 397
rect 399 396 400 397
rect 400 396 401 397
rect 401 396 402 397
rect 402 396 403 397
rect 403 396 404 397
rect 404 396 405 397
rect 405 396 406 397
rect 406 396 407 397
rect 407 396 408 397
rect 408 396 409 397
rect 409 396 410 397
rect 410 396 411 397
rect 411 396 412 397
rect 412 396 413 397
rect 413 396 414 397
rect 414 396 415 397
rect 415 396 416 397
rect 416 396 417 397
rect 417 396 418 397
rect 418 396 419 397
rect 419 396 420 397
rect 420 396 421 397
rect 421 396 422 397
rect 422 396 423 397
rect 423 396 424 397
rect 424 396 425 397
rect 425 396 426 397
rect 426 396 427 397
rect 427 396 428 397
rect 428 396 429 397
rect 429 396 430 397
rect 430 396 431 397
rect 431 396 432 397
rect 432 396 433 397
rect 433 396 434 397
rect 434 396 435 397
rect 435 396 436 397
rect 436 396 437 397
rect 437 396 438 397
rect 438 396 439 397
rect 439 396 440 397
rect 440 396 441 397
rect 441 396 442 397
rect 442 396 443 397
rect 443 396 444 397
rect 444 396 445 397
rect 445 396 446 397
rect 446 396 447 397
rect 447 396 448 397
rect 448 396 449 397
rect 449 396 450 397
rect 450 396 451 397
rect 451 396 452 397
rect 452 396 453 397
rect 453 396 454 397
rect 454 396 455 397
rect 455 396 456 397
rect 456 396 457 397
rect 457 396 458 397
rect 458 396 459 397
rect 459 396 460 397
rect 460 396 461 397
rect 461 396 462 397
rect 462 396 463 397
rect 463 396 464 397
rect 464 396 465 397
rect 465 396 466 397
rect 466 396 467 397
rect 467 396 468 397
rect 468 396 469 397
rect 469 396 470 397
rect 470 396 471 397
rect 471 396 472 397
rect 472 396 473 397
rect 473 396 474 397
rect 474 396 475 397
rect 476 396 477 397
rect 477 396 478 397
rect 478 396 479 397
rect 115 395 116 396
rect 116 395 117 396
rect 117 395 118 396
rect 118 395 119 396
rect 119 395 120 396
rect 120 395 121 396
rect 121 395 122 396
rect 122 395 123 396
rect 123 395 124 396
rect 124 395 125 396
rect 125 395 126 396
rect 126 395 127 396
rect 127 395 128 396
rect 128 395 129 396
rect 173 395 174 396
rect 174 395 175 396
rect 175 395 176 396
rect 176 395 177 396
rect 177 395 178 396
rect 178 395 179 396
rect 179 395 180 396
rect 180 395 181 396
rect 181 395 182 396
rect 182 395 183 396
rect 183 395 184 396
rect 184 395 185 396
rect 185 395 186 396
rect 186 395 187 396
rect 187 395 188 396
rect 188 395 189 396
rect 341 395 342 396
rect 342 395 343 396
rect 343 395 344 396
rect 344 395 345 396
rect 345 395 346 396
rect 346 395 347 396
rect 347 395 348 396
rect 348 395 349 396
rect 349 395 350 396
rect 350 395 351 396
rect 351 395 352 396
rect 353 395 354 396
rect 354 395 355 396
rect 355 395 356 396
rect 356 395 357 396
rect 357 395 358 396
rect 358 395 359 396
rect 359 395 360 396
rect 360 395 361 396
rect 361 395 362 396
rect 362 395 363 396
rect 363 395 364 396
rect 364 395 365 396
rect 365 395 366 396
rect 366 395 367 396
rect 367 395 368 396
rect 368 395 369 396
rect 384 395 385 396
rect 385 395 386 396
rect 386 395 387 396
rect 387 395 388 396
rect 388 395 389 396
rect 389 395 390 396
rect 390 395 391 396
rect 391 395 392 396
rect 392 395 393 396
rect 393 395 394 396
rect 394 395 395 396
rect 395 395 396 396
rect 396 395 397 396
rect 397 395 398 396
rect 398 395 399 396
rect 399 395 400 396
rect 400 395 401 396
rect 401 395 402 396
rect 402 395 403 396
rect 403 395 404 396
rect 404 395 405 396
rect 405 395 406 396
rect 406 395 407 396
rect 407 395 408 396
rect 408 395 409 396
rect 409 395 410 396
rect 410 395 411 396
rect 411 395 412 396
rect 412 395 413 396
rect 413 395 414 396
rect 414 395 415 396
rect 415 395 416 396
rect 416 395 417 396
rect 417 395 418 396
rect 418 395 419 396
rect 419 395 420 396
rect 420 395 421 396
rect 421 395 422 396
rect 422 395 423 396
rect 423 395 424 396
rect 424 395 425 396
rect 425 395 426 396
rect 426 395 427 396
rect 427 395 428 396
rect 428 395 429 396
rect 429 395 430 396
rect 430 395 431 396
rect 431 395 432 396
rect 432 395 433 396
rect 433 395 434 396
rect 434 395 435 396
rect 435 395 436 396
rect 436 395 437 396
rect 437 395 438 396
rect 438 395 439 396
rect 439 395 440 396
rect 440 395 441 396
rect 441 395 442 396
rect 442 395 443 396
rect 443 395 444 396
rect 444 395 445 396
rect 445 395 446 396
rect 446 395 447 396
rect 447 395 448 396
rect 448 395 449 396
rect 449 395 450 396
rect 450 395 451 396
rect 451 395 452 396
rect 452 395 453 396
rect 453 395 454 396
rect 454 395 455 396
rect 455 395 456 396
rect 456 395 457 396
rect 457 395 458 396
rect 458 395 459 396
rect 459 395 460 396
rect 460 395 461 396
rect 461 395 462 396
rect 462 395 463 396
rect 463 395 464 396
rect 464 395 465 396
rect 465 395 466 396
rect 466 395 467 396
rect 467 395 468 396
rect 468 395 469 396
rect 469 395 470 396
rect 470 395 471 396
rect 471 395 472 396
rect 472 395 473 396
rect 473 395 474 396
rect 474 395 475 396
rect 475 395 476 396
rect 476 395 477 396
rect 477 395 478 396
rect 478 395 479 396
rect 479 395 480 396
rect 480 395 481 396
rect 481 395 482 396
rect 482 395 483 396
rect 483 395 484 396
rect 484 395 485 396
rect 485 395 486 396
rect 486 395 487 396
rect 487 395 488 396
rect 115 394 116 395
rect 116 394 117 395
rect 117 394 118 395
rect 118 394 119 395
rect 119 394 120 395
rect 120 394 121 395
rect 121 394 122 395
rect 122 394 123 395
rect 123 394 124 395
rect 124 394 125 395
rect 173 394 174 395
rect 174 394 175 395
rect 175 394 176 395
rect 176 394 177 395
rect 177 394 178 395
rect 178 394 179 395
rect 179 394 180 395
rect 180 394 181 395
rect 181 394 182 395
rect 182 394 183 395
rect 183 394 184 395
rect 184 394 185 395
rect 185 394 186 395
rect 186 394 187 395
rect 341 394 342 395
rect 342 394 343 395
rect 343 394 344 395
rect 344 394 345 395
rect 345 394 346 395
rect 346 394 347 395
rect 347 394 348 395
rect 348 394 349 395
rect 349 394 350 395
rect 350 394 351 395
rect 351 394 352 395
rect 353 394 354 395
rect 354 394 355 395
rect 355 394 356 395
rect 356 394 357 395
rect 357 394 358 395
rect 358 394 359 395
rect 359 394 360 395
rect 360 394 361 395
rect 361 394 362 395
rect 362 394 363 395
rect 363 394 364 395
rect 364 394 365 395
rect 365 394 366 395
rect 366 394 367 395
rect 367 394 368 395
rect 368 394 369 395
rect 384 394 385 395
rect 385 394 386 395
rect 386 394 387 395
rect 387 394 388 395
rect 388 394 389 395
rect 389 394 390 395
rect 390 394 391 395
rect 391 394 392 395
rect 392 394 393 395
rect 393 394 394 395
rect 394 394 395 395
rect 395 394 396 395
rect 396 394 397 395
rect 397 394 398 395
rect 398 394 399 395
rect 399 394 400 395
rect 400 394 401 395
rect 401 394 402 395
rect 402 394 403 395
rect 403 394 404 395
rect 404 394 405 395
rect 405 394 406 395
rect 406 394 407 395
rect 407 394 408 395
rect 408 394 409 395
rect 409 394 410 395
rect 410 394 411 395
rect 411 394 412 395
rect 412 394 413 395
rect 413 394 414 395
rect 414 394 415 395
rect 415 394 416 395
rect 416 394 417 395
rect 417 394 418 395
rect 418 394 419 395
rect 419 394 420 395
rect 420 394 421 395
rect 421 394 422 395
rect 422 394 423 395
rect 423 394 424 395
rect 424 394 425 395
rect 425 394 426 395
rect 426 394 427 395
rect 427 394 428 395
rect 428 394 429 395
rect 429 394 430 395
rect 430 394 431 395
rect 431 394 432 395
rect 432 394 433 395
rect 433 394 434 395
rect 434 394 435 395
rect 435 394 436 395
rect 436 394 437 395
rect 437 394 438 395
rect 438 394 439 395
rect 439 394 440 395
rect 440 394 441 395
rect 441 394 442 395
rect 442 394 443 395
rect 443 394 444 395
rect 444 394 445 395
rect 445 394 446 395
rect 446 394 447 395
rect 447 394 448 395
rect 448 394 449 395
rect 449 394 450 395
rect 450 394 451 395
rect 451 394 452 395
rect 452 394 453 395
rect 453 394 454 395
rect 454 394 455 395
rect 455 394 456 395
rect 456 394 457 395
rect 457 394 458 395
rect 458 394 459 395
rect 459 394 460 395
rect 460 394 461 395
rect 461 394 462 395
rect 462 394 463 395
rect 463 394 464 395
rect 464 394 465 395
rect 465 394 466 395
rect 466 394 467 395
rect 467 394 468 395
rect 468 394 469 395
rect 469 394 470 395
rect 470 394 471 395
rect 471 394 472 395
rect 472 394 473 395
rect 473 394 474 395
rect 474 394 475 395
rect 475 394 476 395
rect 476 394 477 395
rect 477 394 478 395
rect 478 394 479 395
rect 479 394 480 395
rect 480 394 481 395
rect 481 394 482 395
rect 482 394 483 395
rect 483 394 484 395
rect 484 394 485 395
rect 485 394 486 395
rect 486 394 487 395
rect 487 394 488 395
rect 111 393 112 394
rect 112 393 113 394
rect 113 393 114 394
rect 114 393 115 394
rect 115 393 116 394
rect 116 393 117 394
rect 117 393 118 394
rect 118 393 119 394
rect 119 393 120 394
rect 120 393 121 394
rect 121 393 122 394
rect 122 393 123 394
rect 123 393 124 394
rect 124 393 125 394
rect 169 393 170 394
rect 170 393 171 394
rect 171 393 172 394
rect 172 393 173 394
rect 173 393 174 394
rect 174 393 175 394
rect 175 393 176 394
rect 176 393 177 394
rect 177 393 178 394
rect 178 393 179 394
rect 179 393 180 394
rect 180 393 181 394
rect 181 393 182 394
rect 182 393 183 394
rect 183 393 184 394
rect 184 393 185 394
rect 185 393 186 394
rect 186 393 187 394
rect 339 393 340 394
rect 340 393 341 394
rect 341 393 342 394
rect 342 393 343 394
rect 343 393 344 394
rect 344 393 345 394
rect 345 393 346 394
rect 346 393 347 394
rect 347 393 348 394
rect 348 393 349 394
rect 349 393 350 394
rect 350 393 351 394
rect 351 393 352 394
rect 353 393 354 394
rect 354 393 355 394
rect 355 393 356 394
rect 356 393 357 394
rect 357 393 358 394
rect 358 393 359 394
rect 359 393 360 394
rect 360 393 361 394
rect 361 393 362 394
rect 362 393 363 394
rect 363 393 364 394
rect 364 393 365 394
rect 365 393 366 394
rect 366 393 367 394
rect 367 393 368 394
rect 368 393 369 394
rect 383 393 384 394
rect 384 393 385 394
rect 385 393 386 394
rect 386 393 387 394
rect 387 393 388 394
rect 388 393 389 394
rect 389 393 390 394
rect 390 393 391 394
rect 391 393 392 394
rect 392 393 393 394
rect 393 393 394 394
rect 394 393 395 394
rect 395 393 396 394
rect 396 393 397 394
rect 397 393 398 394
rect 398 393 399 394
rect 399 393 400 394
rect 400 393 401 394
rect 401 393 402 394
rect 402 393 403 394
rect 403 393 404 394
rect 404 393 405 394
rect 405 393 406 394
rect 406 393 407 394
rect 407 393 408 394
rect 408 393 409 394
rect 409 393 410 394
rect 410 393 411 394
rect 411 393 412 394
rect 412 393 413 394
rect 413 393 414 394
rect 414 393 415 394
rect 415 393 416 394
rect 416 393 417 394
rect 417 393 418 394
rect 418 393 419 394
rect 419 393 420 394
rect 420 393 421 394
rect 421 393 422 394
rect 422 393 423 394
rect 423 393 424 394
rect 424 393 425 394
rect 425 393 426 394
rect 426 393 427 394
rect 427 393 428 394
rect 428 393 429 394
rect 429 393 430 394
rect 430 393 431 394
rect 431 393 432 394
rect 432 393 433 394
rect 433 393 434 394
rect 434 393 435 394
rect 435 393 436 394
rect 436 393 437 394
rect 437 393 438 394
rect 438 393 439 394
rect 439 393 440 394
rect 440 393 441 394
rect 441 393 442 394
rect 442 393 443 394
rect 443 393 444 394
rect 444 393 445 394
rect 445 393 446 394
rect 446 393 447 394
rect 447 393 448 394
rect 448 393 449 394
rect 449 393 450 394
rect 450 393 451 394
rect 451 393 452 394
rect 452 393 453 394
rect 453 393 454 394
rect 454 393 455 394
rect 455 393 456 394
rect 456 393 457 394
rect 457 393 458 394
rect 458 393 459 394
rect 459 393 460 394
rect 460 393 461 394
rect 461 393 462 394
rect 462 393 463 394
rect 463 393 464 394
rect 464 393 465 394
rect 465 393 466 394
rect 466 393 467 394
rect 467 393 468 394
rect 468 393 469 394
rect 469 393 470 394
rect 470 393 471 394
rect 471 393 472 394
rect 472 393 473 394
rect 473 393 474 394
rect 474 393 475 394
rect 475 393 476 394
rect 476 393 477 394
rect 477 393 478 394
rect 478 393 479 394
rect 479 393 480 394
rect 480 393 481 394
rect 481 393 482 394
rect 482 393 483 394
rect 483 393 484 394
rect 484 393 485 394
rect 485 393 486 394
rect 486 393 487 394
rect 487 393 488 394
rect 488 393 489 394
rect 489 393 490 394
rect 490 393 491 394
rect 491 393 492 394
rect 492 393 493 394
rect 493 393 494 394
rect 111 392 112 393
rect 112 392 113 393
rect 113 392 114 393
rect 114 392 115 393
rect 115 392 116 393
rect 116 392 117 393
rect 117 392 118 393
rect 118 392 119 393
rect 119 392 120 393
rect 120 392 121 393
rect 121 392 122 393
rect 122 392 123 393
rect 169 392 170 393
rect 170 392 171 393
rect 171 392 172 393
rect 172 392 173 393
rect 173 392 174 393
rect 174 392 175 393
rect 175 392 176 393
rect 176 392 177 393
rect 177 392 178 393
rect 178 392 179 393
rect 179 392 180 393
rect 180 392 181 393
rect 181 392 182 393
rect 182 392 183 393
rect 183 392 184 393
rect 184 392 185 393
rect 339 392 340 393
rect 340 392 341 393
rect 341 392 342 393
rect 342 392 343 393
rect 343 392 344 393
rect 344 392 345 393
rect 345 392 346 393
rect 346 392 347 393
rect 347 392 348 393
rect 348 392 349 393
rect 349 392 350 393
rect 350 392 351 393
rect 351 392 352 393
rect 353 392 354 393
rect 354 392 355 393
rect 355 392 356 393
rect 356 392 357 393
rect 357 392 358 393
rect 358 392 359 393
rect 359 392 360 393
rect 360 392 361 393
rect 361 392 362 393
rect 362 392 363 393
rect 363 392 364 393
rect 364 392 365 393
rect 365 392 366 393
rect 366 392 367 393
rect 383 392 384 393
rect 384 392 385 393
rect 385 392 386 393
rect 386 392 387 393
rect 387 392 388 393
rect 388 392 389 393
rect 389 392 390 393
rect 390 392 391 393
rect 391 392 392 393
rect 392 392 393 393
rect 393 392 394 393
rect 394 392 395 393
rect 395 392 396 393
rect 396 392 397 393
rect 397 392 398 393
rect 398 392 399 393
rect 399 392 400 393
rect 400 392 401 393
rect 401 392 402 393
rect 402 392 403 393
rect 403 392 404 393
rect 404 392 405 393
rect 405 392 406 393
rect 406 392 407 393
rect 407 392 408 393
rect 408 392 409 393
rect 409 392 410 393
rect 410 392 411 393
rect 411 392 412 393
rect 412 392 413 393
rect 413 392 414 393
rect 414 392 415 393
rect 415 392 416 393
rect 416 392 417 393
rect 417 392 418 393
rect 418 392 419 393
rect 419 392 420 393
rect 420 392 421 393
rect 421 392 422 393
rect 422 392 423 393
rect 423 392 424 393
rect 424 392 425 393
rect 425 392 426 393
rect 426 392 427 393
rect 427 392 428 393
rect 428 392 429 393
rect 429 392 430 393
rect 430 392 431 393
rect 431 392 432 393
rect 432 392 433 393
rect 433 392 434 393
rect 434 392 435 393
rect 435 392 436 393
rect 436 392 437 393
rect 437 392 438 393
rect 438 392 439 393
rect 439 392 440 393
rect 441 392 442 393
rect 442 392 443 393
rect 457 392 458 393
rect 458 392 459 393
rect 459 392 460 393
rect 460 392 461 393
rect 461 392 462 393
rect 462 392 463 393
rect 463 392 464 393
rect 464 392 465 393
rect 465 392 466 393
rect 466 392 467 393
rect 467 392 468 393
rect 468 392 469 393
rect 469 392 470 393
rect 470 392 471 393
rect 471 392 472 393
rect 472 392 473 393
rect 473 392 474 393
rect 474 392 475 393
rect 475 392 476 393
rect 476 392 477 393
rect 477 392 478 393
rect 478 392 479 393
rect 479 392 480 393
rect 480 392 481 393
rect 481 392 482 393
rect 482 392 483 393
rect 483 392 484 393
rect 484 392 485 393
rect 485 392 486 393
rect 486 392 487 393
rect 487 392 488 393
rect 488 392 489 393
rect 489 392 490 393
rect 490 392 491 393
rect 491 392 492 393
rect 492 392 493 393
rect 493 392 494 393
rect 109 391 110 392
rect 110 391 111 392
rect 111 391 112 392
rect 112 391 113 392
rect 113 391 114 392
rect 114 391 115 392
rect 115 391 116 392
rect 116 391 117 392
rect 117 391 118 392
rect 118 391 119 392
rect 119 391 120 392
rect 120 391 121 392
rect 121 391 122 392
rect 122 391 123 392
rect 167 391 168 392
rect 168 391 169 392
rect 169 391 170 392
rect 170 391 171 392
rect 171 391 172 392
rect 172 391 173 392
rect 173 391 174 392
rect 174 391 175 392
rect 175 391 176 392
rect 176 391 177 392
rect 177 391 178 392
rect 178 391 179 392
rect 179 391 180 392
rect 180 391 181 392
rect 181 391 182 392
rect 182 391 183 392
rect 183 391 184 392
rect 184 391 185 392
rect 339 391 340 392
rect 340 391 341 392
rect 341 391 342 392
rect 342 391 343 392
rect 343 391 344 392
rect 344 391 345 392
rect 345 391 346 392
rect 346 391 347 392
rect 347 391 348 392
rect 348 391 349 392
rect 349 391 350 392
rect 350 391 351 392
rect 351 391 352 392
rect 353 391 354 392
rect 354 391 355 392
rect 355 391 356 392
rect 356 391 357 392
rect 357 391 358 392
rect 358 391 359 392
rect 359 391 360 392
rect 360 391 361 392
rect 361 391 362 392
rect 362 391 363 392
rect 363 391 364 392
rect 364 391 365 392
rect 365 391 366 392
rect 366 391 367 392
rect 367 391 368 392
rect 368 391 369 392
rect 379 391 380 392
rect 380 391 381 392
rect 381 391 382 392
rect 382 391 383 392
rect 383 391 384 392
rect 384 391 385 392
rect 385 391 386 392
rect 386 391 387 392
rect 387 391 388 392
rect 388 391 389 392
rect 389 391 390 392
rect 390 391 391 392
rect 391 391 392 392
rect 392 391 393 392
rect 393 391 394 392
rect 394 391 395 392
rect 395 391 396 392
rect 396 391 397 392
rect 397 391 398 392
rect 398 391 399 392
rect 399 391 400 392
rect 400 391 401 392
rect 401 391 402 392
rect 402 391 403 392
rect 403 391 404 392
rect 404 391 405 392
rect 405 391 406 392
rect 406 391 407 392
rect 407 391 408 392
rect 408 391 409 392
rect 409 391 410 392
rect 410 391 411 392
rect 411 391 412 392
rect 412 391 413 392
rect 413 391 414 392
rect 414 391 415 392
rect 415 391 416 392
rect 416 391 417 392
rect 417 391 418 392
rect 418 391 419 392
rect 419 391 420 392
rect 420 391 421 392
rect 421 391 422 392
rect 422 391 423 392
rect 423 391 424 392
rect 424 391 425 392
rect 425 391 426 392
rect 426 391 427 392
rect 427 391 428 392
rect 428 391 429 392
rect 429 391 430 392
rect 430 391 431 392
rect 431 391 432 392
rect 432 391 433 392
rect 433 391 434 392
rect 434 391 435 392
rect 435 391 436 392
rect 436 391 437 392
rect 437 391 438 392
rect 438 391 439 392
rect 439 391 440 392
rect 441 391 442 392
rect 442 391 443 392
rect 457 391 458 392
rect 458 391 459 392
rect 459 391 460 392
rect 460 391 461 392
rect 461 391 462 392
rect 462 391 463 392
rect 463 391 464 392
rect 464 391 465 392
rect 465 391 466 392
rect 466 391 467 392
rect 467 391 468 392
rect 468 391 469 392
rect 469 391 470 392
rect 470 391 471 392
rect 471 391 472 392
rect 472 391 473 392
rect 473 391 474 392
rect 474 391 475 392
rect 475 391 476 392
rect 476 391 477 392
rect 477 391 478 392
rect 478 391 479 392
rect 479 391 480 392
rect 480 391 481 392
rect 481 391 482 392
rect 482 391 483 392
rect 483 391 484 392
rect 484 391 485 392
rect 485 391 486 392
rect 486 391 487 392
rect 487 391 488 392
rect 488 391 489 392
rect 489 391 490 392
rect 490 391 491 392
rect 491 391 492 392
rect 492 391 493 392
rect 493 391 494 392
rect 494 391 495 392
rect 495 391 496 392
rect 496 391 497 392
rect 497 391 498 392
rect 498 391 499 392
rect 499 391 500 392
rect 109 390 110 391
rect 110 390 111 391
rect 111 390 112 391
rect 112 390 113 391
rect 113 390 114 391
rect 114 390 115 391
rect 115 390 116 391
rect 116 390 117 391
rect 117 390 118 391
rect 118 390 119 391
rect 119 390 120 391
rect 120 390 121 391
rect 167 390 168 391
rect 168 390 169 391
rect 169 390 170 391
rect 170 390 171 391
rect 171 390 172 391
rect 172 390 173 391
rect 173 390 174 391
rect 174 390 175 391
rect 175 390 176 391
rect 176 390 177 391
rect 177 390 178 391
rect 178 390 179 391
rect 179 390 180 391
rect 180 390 181 391
rect 181 390 182 391
rect 182 390 183 391
rect 339 390 340 391
rect 340 390 341 391
rect 341 390 342 391
rect 342 390 343 391
rect 343 390 344 391
rect 344 390 345 391
rect 345 390 346 391
rect 346 390 347 391
rect 347 390 348 391
rect 348 390 349 391
rect 349 390 350 391
rect 350 390 351 391
rect 351 390 352 391
rect 353 390 354 391
rect 354 390 355 391
rect 355 390 356 391
rect 356 390 357 391
rect 357 390 358 391
rect 358 390 359 391
rect 359 390 360 391
rect 360 390 361 391
rect 361 390 362 391
rect 362 390 363 391
rect 363 390 364 391
rect 364 390 365 391
rect 365 390 366 391
rect 366 390 367 391
rect 367 390 368 391
rect 368 390 369 391
rect 379 390 380 391
rect 380 390 381 391
rect 381 390 382 391
rect 382 390 383 391
rect 383 390 384 391
rect 384 390 385 391
rect 385 390 386 391
rect 386 390 387 391
rect 387 390 388 391
rect 388 390 389 391
rect 389 390 390 391
rect 390 390 391 391
rect 391 390 392 391
rect 392 390 393 391
rect 393 390 394 391
rect 394 390 395 391
rect 395 390 396 391
rect 396 390 397 391
rect 397 390 398 391
rect 398 390 399 391
rect 399 390 400 391
rect 400 390 401 391
rect 401 390 402 391
rect 402 390 403 391
rect 403 390 404 391
rect 404 390 405 391
rect 405 390 406 391
rect 406 390 407 391
rect 407 390 408 391
rect 408 390 409 391
rect 409 390 410 391
rect 410 390 411 391
rect 411 390 412 391
rect 412 390 413 391
rect 413 390 414 391
rect 414 390 415 391
rect 415 390 416 391
rect 416 390 417 391
rect 417 390 418 391
rect 418 390 419 391
rect 419 390 420 391
rect 420 390 421 391
rect 421 390 422 391
rect 422 390 423 391
rect 423 390 424 391
rect 424 390 425 391
rect 425 390 426 391
rect 426 390 427 391
rect 427 390 428 391
rect 465 390 466 391
rect 466 390 467 391
rect 467 390 468 391
rect 468 390 469 391
rect 469 390 470 391
rect 470 390 471 391
rect 471 390 472 391
rect 472 390 473 391
rect 473 390 474 391
rect 474 390 475 391
rect 475 390 476 391
rect 476 390 477 391
rect 477 390 478 391
rect 478 390 479 391
rect 479 390 480 391
rect 480 390 481 391
rect 481 390 482 391
rect 482 390 483 391
rect 483 390 484 391
rect 484 390 485 391
rect 485 390 486 391
rect 486 390 487 391
rect 487 390 488 391
rect 488 390 489 391
rect 489 390 490 391
rect 490 390 491 391
rect 491 390 492 391
rect 492 390 493 391
rect 493 390 494 391
rect 494 390 495 391
rect 495 390 496 391
rect 496 390 497 391
rect 497 390 498 391
rect 498 390 499 391
rect 499 390 500 391
rect 103 389 104 390
rect 104 389 105 390
rect 105 389 106 390
rect 106 389 107 390
rect 107 389 108 390
rect 108 389 109 390
rect 109 389 110 390
rect 110 389 111 390
rect 111 389 112 390
rect 112 389 113 390
rect 113 389 114 390
rect 114 389 115 390
rect 115 389 116 390
rect 116 389 117 390
rect 117 389 118 390
rect 118 389 119 390
rect 119 389 120 390
rect 120 389 121 390
rect 165 389 166 390
rect 166 389 167 390
rect 167 389 168 390
rect 168 389 169 390
rect 169 389 170 390
rect 170 389 171 390
rect 171 389 172 390
rect 172 389 173 390
rect 173 389 174 390
rect 174 389 175 390
rect 175 389 176 390
rect 176 389 177 390
rect 177 389 178 390
rect 178 389 179 390
rect 179 389 180 390
rect 180 389 181 390
rect 181 389 182 390
rect 182 389 183 390
rect 339 389 340 390
rect 340 389 341 390
rect 341 389 342 390
rect 342 389 343 390
rect 343 389 344 390
rect 344 389 345 390
rect 345 389 346 390
rect 346 389 347 390
rect 347 389 348 390
rect 348 389 349 390
rect 349 389 350 390
rect 350 389 351 390
rect 351 389 352 390
rect 353 389 354 390
rect 354 389 355 390
rect 355 389 356 390
rect 356 389 357 390
rect 357 389 358 390
rect 358 389 359 390
rect 359 389 360 390
rect 360 389 361 390
rect 361 389 362 390
rect 362 389 363 390
rect 363 389 364 390
rect 364 389 365 390
rect 365 389 366 390
rect 366 389 367 390
rect 367 389 368 390
rect 368 389 369 390
rect 377 389 378 390
rect 378 389 379 390
rect 379 389 380 390
rect 380 389 381 390
rect 381 389 382 390
rect 382 389 383 390
rect 383 389 384 390
rect 384 389 385 390
rect 385 389 386 390
rect 386 389 387 390
rect 387 389 388 390
rect 388 389 389 390
rect 389 389 390 390
rect 390 389 391 390
rect 391 389 392 390
rect 392 389 393 390
rect 393 389 394 390
rect 394 389 395 390
rect 395 389 396 390
rect 396 389 397 390
rect 397 389 398 390
rect 398 389 399 390
rect 399 389 400 390
rect 400 389 401 390
rect 401 389 402 390
rect 402 389 403 390
rect 403 389 404 390
rect 404 389 405 390
rect 405 389 406 390
rect 406 389 407 390
rect 407 389 408 390
rect 408 389 409 390
rect 409 389 410 390
rect 410 389 411 390
rect 411 389 412 390
rect 412 389 413 390
rect 413 389 414 390
rect 414 389 415 390
rect 415 389 416 390
rect 416 389 417 390
rect 417 389 418 390
rect 418 389 419 390
rect 419 389 420 390
rect 420 389 421 390
rect 421 389 422 390
rect 422 389 423 390
rect 423 389 424 390
rect 424 389 425 390
rect 425 389 426 390
rect 426 389 427 390
rect 427 389 428 390
rect 465 389 466 390
rect 466 389 467 390
rect 467 389 468 390
rect 468 389 469 390
rect 469 389 470 390
rect 470 389 471 390
rect 471 389 472 390
rect 472 389 473 390
rect 473 389 474 390
rect 474 389 475 390
rect 475 389 476 390
rect 476 389 477 390
rect 477 389 478 390
rect 478 389 479 390
rect 479 389 480 390
rect 480 389 481 390
rect 481 389 482 390
rect 482 389 483 390
rect 483 389 484 390
rect 484 389 485 390
rect 485 389 486 390
rect 486 389 487 390
rect 487 389 488 390
rect 488 389 489 390
rect 489 389 490 390
rect 490 389 491 390
rect 491 389 492 390
rect 492 389 493 390
rect 493 389 494 390
rect 494 389 495 390
rect 495 389 496 390
rect 496 389 497 390
rect 497 389 498 390
rect 498 389 499 390
rect 499 389 500 390
rect 500 389 501 390
rect 501 389 502 390
rect 502 389 503 390
rect 103 388 104 389
rect 104 388 105 389
rect 105 388 106 389
rect 106 388 107 389
rect 107 388 108 389
rect 108 388 109 389
rect 109 388 110 389
rect 110 388 111 389
rect 111 388 112 389
rect 112 388 113 389
rect 113 388 114 389
rect 114 388 115 389
rect 115 388 116 389
rect 116 388 117 389
rect 117 388 118 389
rect 165 388 166 389
rect 166 388 167 389
rect 167 388 168 389
rect 168 388 169 389
rect 169 388 170 389
rect 170 388 171 389
rect 171 388 172 389
rect 172 388 173 389
rect 173 388 174 389
rect 174 388 175 389
rect 175 388 176 389
rect 176 388 177 389
rect 177 388 178 389
rect 178 388 179 389
rect 179 388 180 389
rect 180 388 181 389
rect 341 388 342 389
rect 342 388 343 389
rect 343 388 344 389
rect 344 388 345 389
rect 345 388 346 389
rect 346 388 347 389
rect 347 388 348 389
rect 348 388 349 389
rect 349 388 350 389
rect 350 388 351 389
rect 351 388 352 389
rect 353 388 354 389
rect 354 388 355 389
rect 355 388 356 389
rect 356 388 357 389
rect 357 388 358 389
rect 358 388 359 389
rect 359 388 360 389
rect 360 388 361 389
rect 361 388 362 389
rect 362 388 363 389
rect 363 388 364 389
rect 364 388 365 389
rect 365 388 366 389
rect 366 388 367 389
rect 367 388 368 389
rect 368 388 369 389
rect 377 388 378 389
rect 378 388 379 389
rect 379 388 380 389
rect 380 388 381 389
rect 381 388 382 389
rect 382 388 383 389
rect 383 388 384 389
rect 384 388 385 389
rect 385 388 386 389
rect 386 388 387 389
rect 387 388 388 389
rect 388 388 389 389
rect 389 388 390 389
rect 390 388 391 389
rect 391 388 392 389
rect 392 388 393 389
rect 393 388 394 389
rect 394 388 395 389
rect 395 388 396 389
rect 396 388 397 389
rect 397 388 398 389
rect 398 388 399 389
rect 399 388 400 389
rect 400 388 401 389
rect 401 388 402 389
rect 402 388 403 389
rect 403 388 404 389
rect 404 388 405 389
rect 405 388 406 389
rect 406 388 407 389
rect 407 388 408 389
rect 408 388 409 389
rect 409 388 410 389
rect 410 388 411 389
rect 411 388 412 389
rect 412 388 413 389
rect 413 388 414 389
rect 414 388 415 389
rect 415 388 416 389
rect 416 388 417 389
rect 417 388 418 389
rect 418 388 419 389
rect 469 388 470 389
rect 470 388 471 389
rect 471 388 472 389
rect 472 388 473 389
rect 473 388 474 389
rect 474 388 475 389
rect 475 388 476 389
rect 476 388 477 389
rect 477 388 478 389
rect 478 388 479 389
rect 479 388 480 389
rect 480 388 481 389
rect 481 388 482 389
rect 482 388 483 389
rect 483 388 484 389
rect 484 388 485 389
rect 485 388 486 389
rect 486 388 487 389
rect 487 388 488 389
rect 488 388 489 389
rect 489 388 490 389
rect 490 388 491 389
rect 491 388 492 389
rect 492 388 493 389
rect 493 388 494 389
rect 494 388 495 389
rect 495 388 496 389
rect 496 388 497 389
rect 497 388 498 389
rect 498 388 499 389
rect 499 388 500 389
rect 500 388 501 389
rect 501 388 502 389
rect 502 388 503 389
rect 100 387 101 388
rect 101 387 102 388
rect 102 387 103 388
rect 103 387 104 388
rect 104 387 105 388
rect 105 387 106 388
rect 106 387 107 388
rect 107 387 108 388
rect 108 387 109 388
rect 109 387 110 388
rect 110 387 111 388
rect 111 387 112 388
rect 112 387 113 388
rect 113 387 114 388
rect 114 387 115 388
rect 115 387 116 388
rect 116 387 117 388
rect 117 387 118 388
rect 163 387 164 388
rect 164 387 165 388
rect 165 387 166 388
rect 166 387 167 388
rect 167 387 168 388
rect 168 387 169 388
rect 169 387 170 388
rect 170 387 171 388
rect 171 387 172 388
rect 172 387 173 388
rect 173 387 174 388
rect 174 387 175 388
rect 175 387 176 388
rect 176 387 177 388
rect 177 387 178 388
rect 178 387 179 388
rect 179 387 180 388
rect 180 387 181 388
rect 339 387 340 388
rect 340 387 341 388
rect 341 387 342 388
rect 342 387 343 388
rect 343 387 344 388
rect 344 387 345 388
rect 345 387 346 388
rect 346 387 347 388
rect 347 387 348 388
rect 348 387 349 388
rect 349 387 350 388
rect 350 387 351 388
rect 351 387 352 388
rect 352 387 353 388
rect 353 387 354 388
rect 354 387 355 388
rect 355 387 356 388
rect 356 387 357 388
rect 357 387 358 388
rect 358 387 359 388
rect 359 387 360 388
rect 360 387 361 388
rect 361 387 362 388
rect 362 387 363 388
rect 363 387 364 388
rect 364 387 365 388
rect 365 387 366 388
rect 366 387 367 388
rect 367 387 368 388
rect 368 387 369 388
rect 373 387 374 388
rect 374 387 375 388
rect 375 387 376 388
rect 376 387 377 388
rect 377 387 378 388
rect 378 387 379 388
rect 379 387 380 388
rect 380 387 381 388
rect 381 387 382 388
rect 382 387 383 388
rect 383 387 384 388
rect 384 387 385 388
rect 385 387 386 388
rect 386 387 387 388
rect 387 387 388 388
rect 388 387 389 388
rect 389 387 390 388
rect 390 387 391 388
rect 391 387 392 388
rect 392 387 393 388
rect 393 387 394 388
rect 394 387 395 388
rect 395 387 396 388
rect 396 387 397 388
rect 397 387 398 388
rect 398 387 399 388
rect 399 387 400 388
rect 400 387 401 388
rect 401 387 402 388
rect 402 387 403 388
rect 403 387 404 388
rect 404 387 405 388
rect 405 387 406 388
rect 406 387 407 388
rect 407 387 408 388
rect 408 387 409 388
rect 409 387 410 388
rect 410 387 411 388
rect 411 387 412 388
rect 412 387 413 388
rect 413 387 414 388
rect 414 387 415 388
rect 415 387 416 388
rect 416 387 417 388
rect 417 387 418 388
rect 418 387 419 388
rect 469 387 470 388
rect 470 387 471 388
rect 471 387 472 388
rect 472 387 473 388
rect 473 387 474 388
rect 474 387 475 388
rect 475 387 476 388
rect 476 387 477 388
rect 477 387 478 388
rect 478 387 479 388
rect 479 387 480 388
rect 480 387 481 388
rect 481 387 482 388
rect 482 387 483 388
rect 483 387 484 388
rect 484 387 485 388
rect 485 387 486 388
rect 486 387 487 388
rect 487 387 488 388
rect 488 387 489 388
rect 489 387 490 388
rect 490 387 491 388
rect 491 387 492 388
rect 492 387 493 388
rect 493 387 494 388
rect 494 387 495 388
rect 495 387 496 388
rect 496 387 497 388
rect 497 387 498 388
rect 498 387 499 388
rect 499 387 500 388
rect 500 387 501 388
rect 501 387 502 388
rect 502 387 503 388
rect 503 387 504 388
rect 504 387 505 388
rect 505 387 506 388
rect 506 387 507 388
rect 100 386 101 387
rect 101 386 102 387
rect 102 386 103 387
rect 103 386 104 387
rect 104 386 105 387
rect 105 386 106 387
rect 106 386 107 387
rect 107 386 108 387
rect 108 386 109 387
rect 109 386 110 387
rect 110 386 111 387
rect 111 386 112 387
rect 112 386 113 387
rect 113 386 114 387
rect 163 386 164 387
rect 164 386 165 387
rect 165 386 166 387
rect 166 386 167 387
rect 167 386 168 387
rect 168 386 169 387
rect 169 386 170 387
rect 170 386 171 387
rect 171 386 172 387
rect 172 386 173 387
rect 173 386 174 387
rect 174 386 175 387
rect 175 386 176 387
rect 176 386 177 387
rect 177 386 178 387
rect 178 386 179 387
rect 339 386 340 387
rect 340 386 341 387
rect 341 386 342 387
rect 342 386 343 387
rect 343 386 344 387
rect 344 386 345 387
rect 345 386 346 387
rect 346 386 347 387
rect 347 386 348 387
rect 348 386 349 387
rect 349 386 350 387
rect 350 386 351 387
rect 351 386 352 387
rect 352 386 353 387
rect 353 386 354 387
rect 354 386 355 387
rect 355 386 356 387
rect 356 386 357 387
rect 357 386 358 387
rect 358 386 359 387
rect 359 386 360 387
rect 360 386 361 387
rect 361 386 362 387
rect 362 386 363 387
rect 363 386 364 387
rect 364 386 365 387
rect 365 386 366 387
rect 366 386 367 387
rect 367 386 368 387
rect 368 386 369 387
rect 373 386 374 387
rect 374 386 375 387
rect 375 386 376 387
rect 376 386 377 387
rect 377 386 378 387
rect 378 386 379 387
rect 379 386 380 387
rect 380 386 381 387
rect 381 386 382 387
rect 382 386 383 387
rect 383 386 384 387
rect 384 386 385 387
rect 385 386 386 387
rect 386 386 387 387
rect 387 386 388 387
rect 388 386 389 387
rect 389 386 390 387
rect 390 386 391 387
rect 391 386 392 387
rect 392 386 393 387
rect 393 386 394 387
rect 394 386 395 387
rect 395 386 396 387
rect 396 386 397 387
rect 397 386 398 387
rect 398 386 399 387
rect 399 386 400 387
rect 400 386 401 387
rect 401 386 402 387
rect 402 386 403 387
rect 403 386 404 387
rect 404 386 405 387
rect 405 386 406 387
rect 406 386 407 387
rect 407 386 408 387
rect 408 386 409 387
rect 409 386 410 387
rect 410 386 411 387
rect 411 386 412 387
rect 474 386 475 387
rect 475 386 476 387
rect 476 386 477 387
rect 477 386 478 387
rect 478 386 479 387
rect 479 386 480 387
rect 480 386 481 387
rect 481 386 482 387
rect 482 386 483 387
rect 483 386 484 387
rect 484 386 485 387
rect 485 386 486 387
rect 486 386 487 387
rect 487 386 488 387
rect 488 386 489 387
rect 489 386 490 387
rect 490 386 491 387
rect 491 386 492 387
rect 492 386 493 387
rect 493 386 494 387
rect 494 386 495 387
rect 495 386 496 387
rect 496 386 497 387
rect 497 386 498 387
rect 498 386 499 387
rect 499 386 500 387
rect 500 386 501 387
rect 501 386 502 387
rect 502 386 503 387
rect 503 386 504 387
rect 504 386 505 387
rect 505 386 506 387
rect 506 386 507 387
rect 98 385 99 386
rect 99 385 100 386
rect 100 385 101 386
rect 101 385 102 386
rect 102 385 103 386
rect 103 385 104 386
rect 104 385 105 386
rect 105 385 106 386
rect 106 385 107 386
rect 107 385 108 386
rect 108 385 109 386
rect 109 385 110 386
rect 110 385 111 386
rect 111 385 112 386
rect 112 385 113 386
rect 113 385 114 386
rect 162 385 163 386
rect 163 385 164 386
rect 164 385 165 386
rect 165 385 166 386
rect 166 385 167 386
rect 167 385 168 386
rect 168 385 169 386
rect 169 385 170 386
rect 170 385 171 386
rect 171 385 172 386
rect 172 385 173 386
rect 173 385 174 386
rect 174 385 175 386
rect 175 385 176 386
rect 176 385 177 386
rect 177 385 178 386
rect 178 385 179 386
rect 339 385 340 386
rect 340 385 341 386
rect 341 385 342 386
rect 342 385 343 386
rect 343 385 344 386
rect 344 385 345 386
rect 345 385 346 386
rect 346 385 347 386
rect 347 385 348 386
rect 348 385 349 386
rect 349 385 350 386
rect 350 385 351 386
rect 351 385 352 386
rect 352 385 353 386
rect 353 385 354 386
rect 354 385 355 386
rect 355 385 356 386
rect 356 385 357 386
rect 357 385 358 386
rect 358 385 359 386
rect 359 385 360 386
rect 360 385 361 386
rect 361 385 362 386
rect 362 385 363 386
rect 363 385 364 386
rect 364 385 365 386
rect 365 385 366 386
rect 366 385 367 386
rect 367 385 368 386
rect 368 385 369 386
rect 369 385 370 386
rect 370 385 371 386
rect 371 385 372 386
rect 372 385 373 386
rect 373 385 374 386
rect 374 385 375 386
rect 375 385 376 386
rect 376 385 377 386
rect 377 385 378 386
rect 378 385 379 386
rect 379 385 380 386
rect 380 385 381 386
rect 381 385 382 386
rect 382 385 383 386
rect 383 385 384 386
rect 384 385 385 386
rect 385 385 386 386
rect 386 385 387 386
rect 387 385 388 386
rect 388 385 389 386
rect 389 385 390 386
rect 390 385 391 386
rect 391 385 392 386
rect 392 385 393 386
rect 393 385 394 386
rect 394 385 395 386
rect 395 385 396 386
rect 396 385 397 386
rect 397 385 398 386
rect 398 385 399 386
rect 399 385 400 386
rect 400 385 401 386
rect 401 385 402 386
rect 402 385 403 386
rect 403 385 404 386
rect 404 385 405 386
rect 405 385 406 386
rect 406 385 407 386
rect 407 385 408 386
rect 408 385 409 386
rect 409 385 410 386
rect 410 385 411 386
rect 411 385 412 386
rect 474 385 475 386
rect 475 385 476 386
rect 476 385 477 386
rect 477 385 478 386
rect 478 385 479 386
rect 479 385 480 386
rect 480 385 481 386
rect 481 385 482 386
rect 482 385 483 386
rect 483 385 484 386
rect 484 385 485 386
rect 485 385 486 386
rect 486 385 487 386
rect 487 385 488 386
rect 488 385 489 386
rect 489 385 490 386
rect 490 385 491 386
rect 491 385 492 386
rect 492 385 493 386
rect 493 385 494 386
rect 494 385 495 386
rect 495 385 496 386
rect 496 385 497 386
rect 497 385 498 386
rect 498 385 499 386
rect 499 385 500 386
rect 500 385 501 386
rect 501 385 502 386
rect 502 385 503 386
rect 503 385 504 386
rect 504 385 505 386
rect 505 385 506 386
rect 506 385 507 386
rect 507 385 508 386
rect 508 385 509 386
rect 98 384 99 385
rect 99 384 100 385
rect 100 384 101 385
rect 101 384 102 385
rect 102 384 103 385
rect 103 384 104 385
rect 104 384 105 385
rect 105 384 106 385
rect 106 384 107 385
rect 107 384 108 385
rect 108 384 109 385
rect 109 384 110 385
rect 110 384 111 385
rect 111 384 112 385
rect 162 384 163 385
rect 163 384 164 385
rect 164 384 165 385
rect 165 384 166 385
rect 166 384 167 385
rect 167 384 168 385
rect 168 384 169 385
rect 169 384 170 385
rect 170 384 171 385
rect 171 384 172 385
rect 172 384 173 385
rect 173 384 174 385
rect 174 384 175 385
rect 175 384 176 385
rect 176 384 177 385
rect 339 384 340 385
rect 340 384 341 385
rect 341 384 342 385
rect 342 384 343 385
rect 343 384 344 385
rect 344 384 345 385
rect 345 384 346 385
rect 346 384 347 385
rect 347 384 348 385
rect 348 384 349 385
rect 349 384 350 385
rect 350 384 351 385
rect 351 384 352 385
rect 352 384 353 385
rect 353 384 354 385
rect 354 384 355 385
rect 355 384 356 385
rect 356 384 357 385
rect 357 384 358 385
rect 358 384 359 385
rect 359 384 360 385
rect 360 384 361 385
rect 361 384 362 385
rect 362 384 363 385
rect 363 384 364 385
rect 364 384 365 385
rect 365 384 366 385
rect 366 384 367 385
rect 367 384 368 385
rect 368 384 369 385
rect 369 384 370 385
rect 370 384 371 385
rect 371 384 372 385
rect 372 384 373 385
rect 373 384 374 385
rect 374 384 375 385
rect 375 384 376 385
rect 376 384 377 385
rect 377 384 378 385
rect 378 384 379 385
rect 379 384 380 385
rect 380 384 381 385
rect 381 384 382 385
rect 382 384 383 385
rect 383 384 384 385
rect 384 384 385 385
rect 385 384 386 385
rect 386 384 387 385
rect 387 384 388 385
rect 388 384 389 385
rect 389 384 390 385
rect 390 384 391 385
rect 391 384 392 385
rect 392 384 393 385
rect 393 384 394 385
rect 394 384 395 385
rect 395 384 396 385
rect 396 384 397 385
rect 397 384 398 385
rect 398 384 399 385
rect 399 384 400 385
rect 400 384 401 385
rect 401 384 402 385
rect 402 384 403 385
rect 403 384 404 385
rect 404 384 405 385
rect 405 384 406 385
rect 476 384 477 385
rect 477 384 478 385
rect 478 384 479 385
rect 479 384 480 385
rect 480 384 481 385
rect 481 384 482 385
rect 482 384 483 385
rect 483 384 484 385
rect 484 384 485 385
rect 485 384 486 385
rect 486 384 487 385
rect 487 384 488 385
rect 488 384 489 385
rect 489 384 490 385
rect 490 384 491 385
rect 491 384 492 385
rect 492 384 493 385
rect 493 384 494 385
rect 494 384 495 385
rect 495 384 496 385
rect 496 384 497 385
rect 497 384 498 385
rect 498 384 499 385
rect 499 384 500 385
rect 500 384 501 385
rect 501 384 502 385
rect 502 384 503 385
rect 503 384 504 385
rect 504 384 505 385
rect 505 384 506 385
rect 506 384 507 385
rect 507 384 508 385
rect 508 384 509 385
rect 92 383 93 384
rect 93 383 94 384
rect 94 383 95 384
rect 95 383 96 384
rect 96 383 97 384
rect 97 383 98 384
rect 98 383 99 384
rect 99 383 100 384
rect 100 383 101 384
rect 101 383 102 384
rect 102 383 103 384
rect 103 383 104 384
rect 104 383 105 384
rect 105 383 106 384
rect 106 383 107 384
rect 107 383 108 384
rect 108 383 109 384
rect 109 383 110 384
rect 110 383 111 384
rect 111 383 112 384
rect 158 383 159 384
rect 159 383 160 384
rect 160 383 161 384
rect 161 383 162 384
rect 162 383 163 384
rect 163 383 164 384
rect 164 383 165 384
rect 165 383 166 384
rect 166 383 167 384
rect 167 383 168 384
rect 168 383 169 384
rect 169 383 170 384
rect 170 383 171 384
rect 171 383 172 384
rect 172 383 173 384
rect 173 383 174 384
rect 174 383 175 384
rect 175 383 176 384
rect 176 383 177 384
rect 339 383 340 384
rect 340 383 341 384
rect 341 383 342 384
rect 342 383 343 384
rect 343 383 344 384
rect 344 383 345 384
rect 345 383 346 384
rect 346 383 347 384
rect 347 383 348 384
rect 348 383 349 384
rect 349 383 350 384
rect 350 383 351 384
rect 351 383 352 384
rect 352 383 353 384
rect 353 383 354 384
rect 354 383 355 384
rect 355 383 356 384
rect 356 383 357 384
rect 357 383 358 384
rect 358 383 359 384
rect 359 383 360 384
rect 360 383 361 384
rect 361 383 362 384
rect 362 383 363 384
rect 363 383 364 384
rect 364 383 365 384
rect 365 383 366 384
rect 366 383 367 384
rect 367 383 368 384
rect 368 383 369 384
rect 369 383 370 384
rect 370 383 371 384
rect 371 383 372 384
rect 372 383 373 384
rect 373 383 374 384
rect 374 383 375 384
rect 375 383 376 384
rect 376 383 377 384
rect 377 383 378 384
rect 378 383 379 384
rect 379 383 380 384
rect 380 383 381 384
rect 381 383 382 384
rect 382 383 383 384
rect 383 383 384 384
rect 384 383 385 384
rect 385 383 386 384
rect 386 383 387 384
rect 387 383 388 384
rect 388 383 389 384
rect 389 383 390 384
rect 390 383 391 384
rect 391 383 392 384
rect 392 383 393 384
rect 393 383 394 384
rect 394 383 395 384
rect 395 383 396 384
rect 396 383 397 384
rect 397 383 398 384
rect 398 383 399 384
rect 399 383 400 384
rect 400 383 401 384
rect 401 383 402 384
rect 402 383 403 384
rect 403 383 404 384
rect 404 383 405 384
rect 405 383 406 384
rect 476 383 477 384
rect 477 383 478 384
rect 478 383 479 384
rect 479 383 480 384
rect 480 383 481 384
rect 481 383 482 384
rect 482 383 483 384
rect 483 383 484 384
rect 484 383 485 384
rect 485 383 486 384
rect 486 383 487 384
rect 487 383 488 384
rect 488 383 489 384
rect 489 383 490 384
rect 490 383 491 384
rect 491 383 492 384
rect 492 383 493 384
rect 493 383 494 384
rect 494 383 495 384
rect 495 383 496 384
rect 496 383 497 384
rect 497 383 498 384
rect 498 383 499 384
rect 499 383 500 384
rect 500 383 501 384
rect 501 383 502 384
rect 502 383 503 384
rect 503 383 504 384
rect 504 383 505 384
rect 505 383 506 384
rect 506 383 507 384
rect 507 383 508 384
rect 508 383 509 384
rect 509 383 510 384
rect 510 383 511 384
rect 511 383 512 384
rect 512 383 513 384
rect 92 382 93 383
rect 93 382 94 383
rect 94 382 95 383
rect 95 382 96 383
rect 96 382 97 383
rect 97 382 98 383
rect 98 382 99 383
rect 99 382 100 383
rect 100 382 101 383
rect 101 382 102 383
rect 102 382 103 383
rect 103 382 104 383
rect 104 382 105 383
rect 105 382 106 383
rect 106 382 107 383
rect 107 382 108 383
rect 158 382 159 383
rect 159 382 160 383
rect 160 382 161 383
rect 161 382 162 383
rect 162 382 163 383
rect 163 382 164 383
rect 164 382 165 383
rect 165 382 166 383
rect 166 382 167 383
rect 167 382 168 383
rect 168 382 169 383
rect 169 382 170 383
rect 170 382 171 383
rect 171 382 172 383
rect 172 382 173 383
rect 173 382 174 383
rect 174 382 175 383
rect 175 382 176 383
rect 339 382 340 383
rect 340 382 341 383
rect 341 382 342 383
rect 342 382 343 383
rect 343 382 344 383
rect 344 382 345 383
rect 345 382 346 383
rect 346 382 347 383
rect 347 382 348 383
rect 348 382 349 383
rect 349 382 350 383
rect 350 382 351 383
rect 351 382 352 383
rect 352 382 353 383
rect 353 382 354 383
rect 354 382 355 383
rect 355 382 356 383
rect 356 382 357 383
rect 357 382 358 383
rect 358 382 359 383
rect 359 382 360 383
rect 360 382 361 383
rect 361 382 362 383
rect 362 382 363 383
rect 363 382 364 383
rect 364 382 365 383
rect 365 382 366 383
rect 366 382 367 383
rect 367 382 368 383
rect 368 382 369 383
rect 369 382 370 383
rect 370 382 371 383
rect 371 382 372 383
rect 372 382 373 383
rect 373 382 374 383
rect 374 382 375 383
rect 375 382 376 383
rect 376 382 377 383
rect 377 382 378 383
rect 378 382 379 383
rect 379 382 380 383
rect 380 382 381 383
rect 381 382 382 383
rect 382 382 383 383
rect 383 382 384 383
rect 384 382 385 383
rect 385 382 386 383
rect 386 382 387 383
rect 387 382 388 383
rect 388 382 389 383
rect 389 382 390 383
rect 390 382 391 383
rect 391 382 392 383
rect 392 382 393 383
rect 393 382 394 383
rect 394 382 395 383
rect 395 382 396 383
rect 396 382 397 383
rect 397 382 398 383
rect 480 382 481 383
rect 481 382 482 383
rect 482 382 483 383
rect 483 382 484 383
rect 484 382 485 383
rect 485 382 486 383
rect 486 382 487 383
rect 487 382 488 383
rect 488 382 489 383
rect 489 382 490 383
rect 490 382 491 383
rect 491 382 492 383
rect 492 382 493 383
rect 493 382 494 383
rect 494 382 495 383
rect 495 382 496 383
rect 496 382 497 383
rect 497 382 498 383
rect 498 382 499 383
rect 499 382 500 383
rect 500 382 501 383
rect 501 382 502 383
rect 502 382 503 383
rect 503 382 504 383
rect 504 382 505 383
rect 505 382 506 383
rect 506 382 507 383
rect 507 382 508 383
rect 508 382 509 383
rect 509 382 510 383
rect 510 382 511 383
rect 511 382 512 383
rect 512 382 513 383
rect 92 381 93 382
rect 93 381 94 382
rect 94 381 95 382
rect 95 381 96 382
rect 96 381 97 382
rect 97 381 98 382
rect 98 381 99 382
rect 99 381 100 382
rect 100 381 101 382
rect 101 381 102 382
rect 102 381 103 382
rect 103 381 104 382
rect 104 381 105 382
rect 105 381 106 382
rect 106 381 107 382
rect 107 381 108 382
rect 158 381 159 382
rect 159 381 160 382
rect 160 381 161 382
rect 161 381 162 382
rect 162 381 163 382
rect 163 381 164 382
rect 164 381 165 382
rect 165 381 166 382
rect 166 381 167 382
rect 167 381 168 382
rect 168 381 169 382
rect 169 381 170 382
rect 170 381 171 382
rect 171 381 172 382
rect 172 381 173 382
rect 173 381 174 382
rect 174 381 175 382
rect 175 381 176 382
rect 339 381 340 382
rect 340 381 341 382
rect 341 381 342 382
rect 342 381 343 382
rect 343 381 344 382
rect 344 381 345 382
rect 345 381 346 382
rect 346 381 347 382
rect 347 381 348 382
rect 348 381 349 382
rect 349 381 350 382
rect 350 381 351 382
rect 351 381 352 382
rect 352 381 353 382
rect 353 381 354 382
rect 354 381 355 382
rect 355 381 356 382
rect 356 381 357 382
rect 357 381 358 382
rect 358 381 359 382
rect 359 381 360 382
rect 360 381 361 382
rect 361 381 362 382
rect 362 381 363 382
rect 363 381 364 382
rect 364 381 365 382
rect 365 381 366 382
rect 366 381 367 382
rect 367 381 368 382
rect 368 381 369 382
rect 369 381 370 382
rect 370 381 371 382
rect 371 381 372 382
rect 372 381 373 382
rect 373 381 374 382
rect 374 381 375 382
rect 375 381 376 382
rect 376 381 377 382
rect 377 381 378 382
rect 378 381 379 382
rect 379 381 380 382
rect 380 381 381 382
rect 381 381 382 382
rect 382 381 383 382
rect 383 381 384 382
rect 384 381 385 382
rect 385 381 386 382
rect 386 381 387 382
rect 387 381 388 382
rect 388 381 389 382
rect 389 381 390 382
rect 390 381 391 382
rect 391 381 392 382
rect 392 381 393 382
rect 393 381 394 382
rect 394 381 395 382
rect 395 381 396 382
rect 396 381 397 382
rect 397 381 398 382
rect 480 381 481 382
rect 481 381 482 382
rect 482 381 483 382
rect 483 381 484 382
rect 484 381 485 382
rect 485 381 486 382
rect 486 381 487 382
rect 487 381 488 382
rect 488 381 489 382
rect 489 381 490 382
rect 490 381 491 382
rect 491 381 492 382
rect 492 381 493 382
rect 493 381 494 382
rect 494 381 495 382
rect 495 381 496 382
rect 496 381 497 382
rect 497 381 498 382
rect 498 381 499 382
rect 499 381 500 382
rect 500 381 501 382
rect 501 381 502 382
rect 502 381 503 382
rect 503 381 504 382
rect 504 381 505 382
rect 505 381 506 382
rect 506 381 507 382
rect 507 381 508 382
rect 508 381 509 382
rect 509 381 510 382
rect 510 381 511 382
rect 511 381 512 382
rect 512 381 513 382
rect 88 380 89 381
rect 89 380 90 381
rect 90 380 91 381
rect 91 380 92 381
rect 92 380 93 381
rect 93 380 94 381
rect 94 380 95 381
rect 95 380 96 381
rect 96 380 97 381
rect 97 380 98 381
rect 98 380 99 381
rect 99 380 100 381
rect 100 380 101 381
rect 101 380 102 381
rect 102 380 103 381
rect 103 380 104 381
rect 104 380 105 381
rect 105 380 106 381
rect 106 380 107 381
rect 107 380 108 381
rect 158 380 159 381
rect 159 380 160 381
rect 160 380 161 381
rect 161 380 162 381
rect 162 380 163 381
rect 163 380 164 381
rect 164 380 165 381
rect 165 380 166 381
rect 166 380 167 381
rect 167 380 168 381
rect 168 380 169 381
rect 169 380 170 381
rect 170 380 171 381
rect 171 380 172 381
rect 172 380 173 381
rect 173 380 174 381
rect 174 380 175 381
rect 175 380 176 381
rect 338 380 339 381
rect 339 380 340 381
rect 340 380 341 381
rect 341 380 342 381
rect 342 380 343 381
rect 343 380 344 381
rect 344 380 345 381
rect 345 380 346 381
rect 346 380 347 381
rect 347 380 348 381
rect 348 380 349 381
rect 349 380 350 381
rect 350 380 351 381
rect 351 380 352 381
rect 352 380 353 381
rect 353 380 354 381
rect 354 380 355 381
rect 355 380 356 381
rect 356 380 357 381
rect 357 380 358 381
rect 358 380 359 381
rect 359 380 360 381
rect 360 380 361 381
rect 361 380 362 381
rect 362 380 363 381
rect 363 380 364 381
rect 364 380 365 381
rect 365 380 366 381
rect 366 380 367 381
rect 367 380 368 381
rect 368 380 369 381
rect 369 380 370 381
rect 370 380 371 381
rect 371 380 372 381
rect 372 380 373 381
rect 373 380 374 381
rect 374 380 375 381
rect 375 380 376 381
rect 376 380 377 381
rect 377 380 378 381
rect 378 380 379 381
rect 379 380 380 381
rect 380 380 381 381
rect 381 380 382 381
rect 382 380 383 381
rect 383 380 384 381
rect 384 380 385 381
rect 385 380 386 381
rect 386 380 387 381
rect 387 380 388 381
rect 388 380 389 381
rect 389 380 390 381
rect 390 380 391 381
rect 391 380 392 381
rect 392 380 393 381
rect 393 380 394 381
rect 394 380 395 381
rect 395 380 396 381
rect 396 380 397 381
rect 397 380 398 381
rect 480 380 481 381
rect 481 380 482 381
rect 482 380 483 381
rect 483 380 484 381
rect 484 380 485 381
rect 485 380 486 381
rect 486 380 487 381
rect 487 380 488 381
rect 488 380 489 381
rect 489 380 490 381
rect 490 380 491 381
rect 491 380 492 381
rect 492 380 493 381
rect 493 380 494 381
rect 494 380 495 381
rect 495 380 496 381
rect 496 380 497 381
rect 497 380 498 381
rect 498 380 499 381
rect 499 380 500 381
rect 500 380 501 381
rect 501 380 502 381
rect 502 380 503 381
rect 503 380 504 381
rect 504 380 505 381
rect 505 380 506 381
rect 506 380 507 381
rect 507 380 508 381
rect 508 380 509 381
rect 509 380 510 381
rect 510 380 511 381
rect 511 380 512 381
rect 512 380 513 381
rect 513 380 514 381
rect 514 380 515 381
rect 88 379 89 380
rect 89 379 90 380
rect 90 379 91 380
rect 91 379 92 380
rect 92 379 93 380
rect 93 379 94 380
rect 94 379 95 380
rect 95 379 96 380
rect 96 379 97 380
rect 97 379 98 380
rect 98 379 99 380
rect 99 379 100 380
rect 100 379 101 380
rect 101 379 102 380
rect 102 379 103 380
rect 103 379 104 380
rect 104 379 105 380
rect 105 379 106 380
rect 158 379 159 380
rect 159 379 160 380
rect 160 379 161 380
rect 161 379 162 380
rect 162 379 163 380
rect 163 379 164 380
rect 164 379 165 380
rect 165 379 166 380
rect 166 379 167 380
rect 167 379 168 380
rect 168 379 169 380
rect 169 379 170 380
rect 170 379 171 380
rect 171 379 172 380
rect 172 379 173 380
rect 173 379 174 380
rect 338 379 339 380
rect 339 379 340 380
rect 340 379 341 380
rect 341 379 342 380
rect 342 379 343 380
rect 343 379 344 380
rect 344 379 345 380
rect 345 379 346 380
rect 346 379 347 380
rect 347 379 348 380
rect 348 379 349 380
rect 349 379 350 380
rect 350 379 351 380
rect 351 379 352 380
rect 352 379 353 380
rect 353 379 354 380
rect 354 379 355 380
rect 355 379 356 380
rect 356 379 357 380
rect 357 379 358 380
rect 358 379 359 380
rect 359 379 360 380
rect 360 379 361 380
rect 361 379 362 380
rect 362 379 363 380
rect 363 379 364 380
rect 364 379 365 380
rect 365 379 366 380
rect 366 379 367 380
rect 367 379 368 380
rect 368 379 369 380
rect 369 379 370 380
rect 370 379 371 380
rect 371 379 372 380
rect 372 379 373 380
rect 373 379 374 380
rect 374 379 375 380
rect 375 379 376 380
rect 376 379 377 380
rect 377 379 378 380
rect 378 379 379 380
rect 379 379 380 380
rect 380 379 381 380
rect 381 379 382 380
rect 382 379 383 380
rect 383 379 384 380
rect 384 379 385 380
rect 385 379 386 380
rect 386 379 387 380
rect 387 379 388 380
rect 388 379 389 380
rect 389 379 390 380
rect 390 379 391 380
rect 391 379 392 380
rect 392 379 393 380
rect 482 379 483 380
rect 483 379 484 380
rect 484 379 485 380
rect 485 379 486 380
rect 486 379 487 380
rect 487 379 488 380
rect 488 379 489 380
rect 489 379 490 380
rect 490 379 491 380
rect 491 379 492 380
rect 492 379 493 380
rect 493 379 494 380
rect 494 379 495 380
rect 495 379 496 380
rect 496 379 497 380
rect 497 379 498 380
rect 498 379 499 380
rect 499 379 500 380
rect 500 379 501 380
rect 501 379 502 380
rect 502 379 503 380
rect 503 379 504 380
rect 504 379 505 380
rect 505 379 506 380
rect 506 379 507 380
rect 507 379 508 380
rect 508 379 509 380
rect 509 379 510 380
rect 510 379 511 380
rect 511 379 512 380
rect 512 379 513 380
rect 513 379 514 380
rect 514 379 515 380
rect 85 378 86 379
rect 86 378 87 379
rect 87 378 88 379
rect 88 378 89 379
rect 89 378 90 379
rect 90 378 91 379
rect 91 378 92 379
rect 92 378 93 379
rect 93 378 94 379
rect 94 378 95 379
rect 95 378 96 379
rect 96 378 97 379
rect 97 378 98 379
rect 98 378 99 379
rect 99 378 100 379
rect 100 378 101 379
rect 101 378 102 379
rect 102 378 103 379
rect 103 378 104 379
rect 104 378 105 379
rect 105 378 106 379
rect 154 378 155 379
rect 155 378 156 379
rect 156 378 157 379
rect 157 378 158 379
rect 158 378 159 379
rect 159 378 160 379
rect 160 378 161 379
rect 161 378 162 379
rect 162 378 163 379
rect 163 378 164 379
rect 164 378 165 379
rect 165 378 166 379
rect 166 378 167 379
rect 167 378 168 379
rect 168 378 169 379
rect 169 378 170 379
rect 170 378 171 379
rect 171 378 172 379
rect 172 378 173 379
rect 173 378 174 379
rect 338 378 339 379
rect 339 378 340 379
rect 340 378 341 379
rect 341 378 342 379
rect 342 378 343 379
rect 343 378 344 379
rect 344 378 345 379
rect 345 378 346 379
rect 346 378 347 379
rect 347 378 348 379
rect 348 378 349 379
rect 349 378 350 379
rect 350 378 351 379
rect 351 378 352 379
rect 352 378 353 379
rect 353 378 354 379
rect 354 378 355 379
rect 355 378 356 379
rect 356 378 357 379
rect 357 378 358 379
rect 358 378 359 379
rect 359 378 360 379
rect 360 378 361 379
rect 361 378 362 379
rect 362 378 363 379
rect 363 378 364 379
rect 364 378 365 379
rect 365 378 366 379
rect 366 378 367 379
rect 367 378 368 379
rect 368 378 369 379
rect 369 378 370 379
rect 370 378 371 379
rect 371 378 372 379
rect 372 378 373 379
rect 373 378 374 379
rect 374 378 375 379
rect 375 378 376 379
rect 376 378 377 379
rect 377 378 378 379
rect 378 378 379 379
rect 379 378 380 379
rect 380 378 381 379
rect 381 378 382 379
rect 382 378 383 379
rect 383 378 384 379
rect 384 378 385 379
rect 385 378 386 379
rect 386 378 387 379
rect 387 378 388 379
rect 388 378 389 379
rect 389 378 390 379
rect 390 378 391 379
rect 391 378 392 379
rect 392 378 393 379
rect 482 378 483 379
rect 483 378 484 379
rect 484 378 485 379
rect 485 378 486 379
rect 486 378 487 379
rect 487 378 488 379
rect 488 378 489 379
rect 489 378 490 379
rect 490 378 491 379
rect 491 378 492 379
rect 492 378 493 379
rect 493 378 494 379
rect 494 378 495 379
rect 495 378 496 379
rect 496 378 497 379
rect 497 378 498 379
rect 498 378 499 379
rect 499 378 500 379
rect 500 378 501 379
rect 501 378 502 379
rect 502 378 503 379
rect 503 378 504 379
rect 504 378 505 379
rect 505 378 506 379
rect 506 378 507 379
rect 507 378 508 379
rect 508 378 509 379
rect 509 378 510 379
rect 510 378 511 379
rect 511 378 512 379
rect 512 378 513 379
rect 513 378 514 379
rect 514 378 515 379
rect 515 378 516 379
rect 85 377 86 378
rect 86 377 87 378
rect 87 377 88 378
rect 88 377 89 378
rect 89 377 90 378
rect 90 377 91 378
rect 91 377 92 378
rect 92 377 93 378
rect 93 377 94 378
rect 94 377 95 378
rect 95 377 96 378
rect 96 377 97 378
rect 97 377 98 378
rect 98 377 99 378
rect 99 377 100 378
rect 100 377 101 378
rect 101 377 102 378
rect 102 377 103 378
rect 154 377 155 378
rect 155 377 156 378
rect 156 377 157 378
rect 157 377 158 378
rect 158 377 159 378
rect 159 377 160 378
rect 160 377 161 378
rect 161 377 162 378
rect 162 377 163 378
rect 163 377 164 378
rect 164 377 165 378
rect 165 377 166 378
rect 166 377 167 378
rect 167 377 168 378
rect 168 377 169 378
rect 169 377 170 378
rect 170 377 171 378
rect 171 377 172 378
rect 338 377 339 378
rect 339 377 340 378
rect 340 377 341 378
rect 341 377 342 378
rect 342 377 343 378
rect 343 377 344 378
rect 344 377 345 378
rect 345 377 346 378
rect 346 377 347 378
rect 347 377 348 378
rect 348 377 349 378
rect 349 377 350 378
rect 350 377 351 378
rect 351 377 352 378
rect 352 377 353 378
rect 353 377 354 378
rect 354 377 355 378
rect 355 377 356 378
rect 356 377 357 378
rect 357 377 358 378
rect 358 377 359 378
rect 359 377 360 378
rect 360 377 361 378
rect 361 377 362 378
rect 362 377 363 378
rect 363 377 364 378
rect 364 377 365 378
rect 365 377 366 378
rect 366 377 367 378
rect 367 377 368 378
rect 368 377 369 378
rect 369 377 370 378
rect 370 377 371 378
rect 371 377 372 378
rect 372 377 373 378
rect 373 377 374 378
rect 374 377 375 378
rect 375 377 376 378
rect 376 377 377 378
rect 377 377 378 378
rect 378 377 379 378
rect 379 377 380 378
rect 380 377 381 378
rect 381 377 382 378
rect 382 377 383 378
rect 383 377 384 378
rect 384 377 385 378
rect 486 377 487 378
rect 487 377 488 378
rect 488 377 489 378
rect 489 377 490 378
rect 490 377 491 378
rect 491 377 492 378
rect 492 377 493 378
rect 493 377 494 378
rect 494 377 495 378
rect 495 377 496 378
rect 496 377 497 378
rect 497 377 498 378
rect 498 377 499 378
rect 499 377 500 378
rect 500 377 501 378
rect 501 377 502 378
rect 502 377 503 378
rect 503 377 504 378
rect 504 377 505 378
rect 505 377 506 378
rect 506 377 507 378
rect 507 377 508 378
rect 508 377 509 378
rect 509 377 510 378
rect 510 377 511 378
rect 511 377 512 378
rect 512 377 513 378
rect 513 377 514 378
rect 514 377 515 378
rect 515 377 516 378
rect 81 376 82 377
rect 82 376 83 377
rect 83 376 84 377
rect 84 376 85 377
rect 85 376 86 377
rect 86 376 87 377
rect 87 376 88 377
rect 88 376 89 377
rect 89 376 90 377
rect 90 376 91 377
rect 91 376 92 377
rect 92 376 93 377
rect 93 376 94 377
rect 94 376 95 377
rect 95 376 96 377
rect 96 376 97 377
rect 97 376 98 377
rect 98 376 99 377
rect 99 376 100 377
rect 100 376 101 377
rect 101 376 102 377
rect 102 376 103 377
rect 152 376 153 377
rect 153 376 154 377
rect 154 376 155 377
rect 155 376 156 377
rect 156 376 157 377
rect 157 376 158 377
rect 158 376 159 377
rect 159 376 160 377
rect 160 376 161 377
rect 161 376 162 377
rect 162 376 163 377
rect 163 376 164 377
rect 164 376 165 377
rect 165 376 166 377
rect 166 376 167 377
rect 167 376 168 377
rect 168 376 169 377
rect 169 376 170 377
rect 170 376 171 377
rect 171 376 172 377
rect 338 376 339 377
rect 339 376 340 377
rect 340 376 341 377
rect 341 376 342 377
rect 342 376 343 377
rect 343 376 344 377
rect 344 376 345 377
rect 345 376 346 377
rect 346 376 347 377
rect 347 376 348 377
rect 348 376 349 377
rect 349 376 350 377
rect 350 376 351 377
rect 351 376 352 377
rect 352 376 353 377
rect 353 376 354 377
rect 354 376 355 377
rect 355 376 356 377
rect 356 376 357 377
rect 357 376 358 377
rect 358 376 359 377
rect 359 376 360 377
rect 360 376 361 377
rect 361 376 362 377
rect 362 376 363 377
rect 363 376 364 377
rect 364 376 365 377
rect 365 376 366 377
rect 366 376 367 377
rect 367 376 368 377
rect 368 376 369 377
rect 369 376 370 377
rect 370 376 371 377
rect 371 376 372 377
rect 372 376 373 377
rect 373 376 374 377
rect 374 376 375 377
rect 375 376 376 377
rect 376 376 377 377
rect 377 376 378 377
rect 378 376 379 377
rect 379 376 380 377
rect 380 376 381 377
rect 381 376 382 377
rect 382 376 383 377
rect 383 376 384 377
rect 384 376 385 377
rect 486 376 487 377
rect 487 376 488 377
rect 488 376 489 377
rect 489 376 490 377
rect 490 376 491 377
rect 491 376 492 377
rect 492 376 493 377
rect 493 376 494 377
rect 494 376 495 377
rect 495 376 496 377
rect 496 376 497 377
rect 497 376 498 377
rect 498 376 499 377
rect 499 376 500 377
rect 500 376 501 377
rect 501 376 502 377
rect 502 376 503 377
rect 503 376 504 377
rect 504 376 505 377
rect 505 376 506 377
rect 506 376 507 377
rect 507 376 508 377
rect 508 376 509 377
rect 509 376 510 377
rect 510 376 511 377
rect 511 376 512 377
rect 512 376 513 377
rect 513 376 514 377
rect 514 376 515 377
rect 515 376 516 377
rect 516 376 517 377
rect 517 376 518 377
rect 81 375 82 376
rect 82 375 83 376
rect 83 375 84 376
rect 84 375 85 376
rect 85 375 86 376
rect 86 375 87 376
rect 87 375 88 376
rect 88 375 89 376
rect 89 375 90 376
rect 90 375 91 376
rect 91 375 92 376
rect 92 375 93 376
rect 93 375 94 376
rect 94 375 95 376
rect 95 375 96 376
rect 96 375 97 376
rect 97 375 98 376
rect 98 375 99 376
rect 152 375 153 376
rect 153 375 154 376
rect 154 375 155 376
rect 155 375 156 376
rect 156 375 157 376
rect 157 375 158 376
rect 158 375 159 376
rect 159 375 160 376
rect 160 375 161 376
rect 161 375 162 376
rect 162 375 163 376
rect 163 375 164 376
rect 164 375 165 376
rect 165 375 166 376
rect 166 375 167 376
rect 167 375 168 376
rect 168 375 169 376
rect 169 375 170 376
rect 338 375 339 376
rect 339 375 340 376
rect 340 375 341 376
rect 341 375 342 376
rect 342 375 343 376
rect 343 375 344 376
rect 344 375 345 376
rect 345 375 346 376
rect 346 375 347 376
rect 347 375 348 376
rect 348 375 349 376
rect 349 375 350 376
rect 350 375 351 376
rect 351 375 352 376
rect 352 375 353 376
rect 353 375 354 376
rect 354 375 355 376
rect 355 375 356 376
rect 356 375 357 376
rect 357 375 358 376
rect 358 375 359 376
rect 359 375 360 376
rect 360 375 361 376
rect 361 375 362 376
rect 362 375 363 376
rect 363 375 364 376
rect 364 375 365 376
rect 365 375 366 376
rect 366 375 367 376
rect 367 375 368 376
rect 368 375 369 376
rect 369 375 370 376
rect 370 375 371 376
rect 371 375 372 376
rect 372 375 373 376
rect 373 375 374 376
rect 374 375 375 376
rect 375 375 376 376
rect 376 375 377 376
rect 377 375 378 376
rect 378 375 379 376
rect 379 375 380 376
rect 487 375 488 376
rect 488 375 489 376
rect 489 375 490 376
rect 490 375 491 376
rect 491 375 492 376
rect 492 375 493 376
rect 493 375 494 376
rect 494 375 495 376
rect 495 375 496 376
rect 496 375 497 376
rect 497 375 498 376
rect 498 375 499 376
rect 499 375 500 376
rect 500 375 501 376
rect 501 375 502 376
rect 502 375 503 376
rect 503 375 504 376
rect 504 375 505 376
rect 505 375 506 376
rect 506 375 507 376
rect 507 375 508 376
rect 508 375 509 376
rect 509 375 510 376
rect 510 375 511 376
rect 511 375 512 376
rect 512 375 513 376
rect 513 375 514 376
rect 514 375 515 376
rect 515 375 516 376
rect 516 375 517 376
rect 517 375 518 376
rect 77 374 78 375
rect 78 374 79 375
rect 79 374 80 375
rect 80 374 81 375
rect 81 374 82 375
rect 82 374 83 375
rect 83 374 84 375
rect 84 374 85 375
rect 85 374 86 375
rect 86 374 87 375
rect 87 374 88 375
rect 88 374 89 375
rect 89 374 90 375
rect 90 374 91 375
rect 91 374 92 375
rect 92 374 93 375
rect 93 374 94 375
rect 94 374 95 375
rect 95 374 96 375
rect 96 374 97 375
rect 97 374 98 375
rect 98 374 99 375
rect 150 374 151 375
rect 151 374 152 375
rect 152 374 153 375
rect 153 374 154 375
rect 154 374 155 375
rect 155 374 156 375
rect 156 374 157 375
rect 157 374 158 375
rect 158 374 159 375
rect 159 374 160 375
rect 160 374 161 375
rect 161 374 162 375
rect 162 374 163 375
rect 163 374 164 375
rect 164 374 165 375
rect 165 374 166 375
rect 166 374 167 375
rect 167 374 168 375
rect 168 374 169 375
rect 169 374 170 375
rect 336 374 337 375
rect 337 374 338 375
rect 338 374 339 375
rect 339 374 340 375
rect 340 374 341 375
rect 341 374 342 375
rect 342 374 343 375
rect 343 374 344 375
rect 344 374 345 375
rect 345 374 346 375
rect 346 374 347 375
rect 347 374 348 375
rect 348 374 349 375
rect 349 374 350 375
rect 350 374 351 375
rect 351 374 352 375
rect 352 374 353 375
rect 353 374 354 375
rect 354 374 355 375
rect 355 374 356 375
rect 356 374 357 375
rect 357 374 358 375
rect 358 374 359 375
rect 359 374 360 375
rect 360 374 361 375
rect 361 374 362 375
rect 362 374 363 375
rect 363 374 364 375
rect 364 374 365 375
rect 365 374 366 375
rect 366 374 367 375
rect 367 374 368 375
rect 368 374 369 375
rect 369 374 370 375
rect 370 374 371 375
rect 371 374 372 375
rect 372 374 373 375
rect 373 374 374 375
rect 374 374 375 375
rect 375 374 376 375
rect 376 374 377 375
rect 377 374 378 375
rect 378 374 379 375
rect 379 374 380 375
rect 487 374 488 375
rect 488 374 489 375
rect 489 374 490 375
rect 490 374 491 375
rect 491 374 492 375
rect 492 374 493 375
rect 493 374 494 375
rect 494 374 495 375
rect 495 374 496 375
rect 496 374 497 375
rect 497 374 498 375
rect 498 374 499 375
rect 499 374 500 375
rect 500 374 501 375
rect 501 374 502 375
rect 502 374 503 375
rect 503 374 504 375
rect 504 374 505 375
rect 505 374 506 375
rect 506 374 507 375
rect 507 374 508 375
rect 508 374 509 375
rect 509 374 510 375
rect 510 374 511 375
rect 511 374 512 375
rect 512 374 513 375
rect 513 374 514 375
rect 514 374 515 375
rect 515 374 516 375
rect 516 374 517 375
rect 517 374 518 375
rect 518 374 519 375
rect 519 374 520 375
rect 77 373 78 374
rect 78 373 79 374
rect 79 373 80 374
rect 80 373 81 374
rect 81 373 82 374
rect 82 373 83 374
rect 83 373 84 374
rect 84 373 85 374
rect 85 373 86 374
rect 86 373 87 374
rect 87 373 88 374
rect 88 373 89 374
rect 89 373 90 374
rect 90 373 91 374
rect 91 373 92 374
rect 92 373 93 374
rect 93 373 94 374
rect 94 373 95 374
rect 150 373 151 374
rect 151 373 152 374
rect 152 373 153 374
rect 153 373 154 374
rect 154 373 155 374
rect 155 373 156 374
rect 156 373 157 374
rect 157 373 158 374
rect 158 373 159 374
rect 159 373 160 374
rect 160 373 161 374
rect 161 373 162 374
rect 162 373 163 374
rect 163 373 164 374
rect 164 373 165 374
rect 165 373 166 374
rect 166 373 167 374
rect 167 373 168 374
rect 336 373 337 374
rect 337 373 338 374
rect 338 373 339 374
rect 339 373 340 374
rect 340 373 341 374
rect 341 373 342 374
rect 342 373 343 374
rect 343 373 344 374
rect 344 373 345 374
rect 345 373 346 374
rect 346 373 347 374
rect 347 373 348 374
rect 348 373 349 374
rect 349 373 350 374
rect 350 373 351 374
rect 351 373 352 374
rect 352 373 353 374
rect 353 373 354 374
rect 354 373 355 374
rect 355 373 356 374
rect 356 373 357 374
rect 357 373 358 374
rect 358 373 359 374
rect 359 373 360 374
rect 360 373 361 374
rect 361 373 362 374
rect 362 373 363 374
rect 363 373 364 374
rect 364 373 365 374
rect 365 373 366 374
rect 366 373 367 374
rect 367 373 368 374
rect 368 373 369 374
rect 369 373 370 374
rect 370 373 371 374
rect 371 373 372 374
rect 489 373 490 374
rect 490 373 491 374
rect 491 373 492 374
rect 492 373 493 374
rect 493 373 494 374
rect 494 373 495 374
rect 495 373 496 374
rect 496 373 497 374
rect 497 373 498 374
rect 498 373 499 374
rect 499 373 500 374
rect 500 373 501 374
rect 501 373 502 374
rect 502 373 503 374
rect 503 373 504 374
rect 504 373 505 374
rect 505 373 506 374
rect 506 373 507 374
rect 507 373 508 374
rect 508 373 509 374
rect 509 373 510 374
rect 510 373 511 374
rect 511 373 512 374
rect 512 373 513 374
rect 513 373 514 374
rect 514 373 515 374
rect 515 373 516 374
rect 516 373 517 374
rect 517 373 518 374
rect 518 373 519 374
rect 519 373 520 374
rect 73 372 74 373
rect 74 372 75 373
rect 75 372 76 373
rect 76 372 77 373
rect 77 372 78 373
rect 78 372 79 373
rect 79 372 80 373
rect 80 372 81 373
rect 81 372 82 373
rect 82 372 83 373
rect 83 372 84 373
rect 84 372 85 373
rect 85 372 86 373
rect 86 372 87 373
rect 87 372 88 373
rect 88 372 89 373
rect 89 372 90 373
rect 90 372 91 373
rect 91 372 92 373
rect 92 372 93 373
rect 93 372 94 373
rect 94 372 95 373
rect 148 372 149 373
rect 149 372 150 373
rect 150 372 151 373
rect 151 372 152 373
rect 152 372 153 373
rect 153 372 154 373
rect 154 372 155 373
rect 155 372 156 373
rect 156 372 157 373
rect 157 372 158 373
rect 158 372 159 373
rect 159 372 160 373
rect 160 372 161 373
rect 161 372 162 373
rect 162 372 163 373
rect 163 372 164 373
rect 164 372 165 373
rect 165 372 166 373
rect 166 372 167 373
rect 167 372 168 373
rect 334 372 335 373
rect 335 372 336 373
rect 336 372 337 373
rect 337 372 338 373
rect 338 372 339 373
rect 339 372 340 373
rect 340 372 341 373
rect 341 372 342 373
rect 342 372 343 373
rect 343 372 344 373
rect 344 372 345 373
rect 345 372 346 373
rect 346 372 347 373
rect 347 372 348 373
rect 348 372 349 373
rect 349 372 350 373
rect 350 372 351 373
rect 351 372 352 373
rect 352 372 353 373
rect 353 372 354 373
rect 354 372 355 373
rect 355 372 356 373
rect 356 372 357 373
rect 357 372 358 373
rect 358 372 359 373
rect 359 372 360 373
rect 360 372 361 373
rect 361 372 362 373
rect 362 372 363 373
rect 363 372 364 373
rect 364 372 365 373
rect 365 372 366 373
rect 366 372 367 373
rect 367 372 368 373
rect 368 372 369 373
rect 369 372 370 373
rect 370 372 371 373
rect 371 372 372 373
rect 489 372 490 373
rect 490 372 491 373
rect 491 372 492 373
rect 492 372 493 373
rect 493 372 494 373
rect 494 372 495 373
rect 495 372 496 373
rect 496 372 497 373
rect 497 372 498 373
rect 498 372 499 373
rect 499 372 500 373
rect 500 372 501 373
rect 501 372 502 373
rect 502 372 503 373
rect 503 372 504 373
rect 504 372 505 373
rect 505 372 506 373
rect 506 372 507 373
rect 507 372 508 373
rect 508 372 509 373
rect 509 372 510 373
rect 510 372 511 373
rect 511 372 512 373
rect 512 372 513 373
rect 513 372 514 373
rect 514 372 515 373
rect 515 372 516 373
rect 516 372 517 373
rect 517 372 518 373
rect 518 372 519 373
rect 519 372 520 373
rect 520 372 521 373
rect 521 372 522 373
rect 73 371 74 372
rect 74 371 75 372
rect 75 371 76 372
rect 76 371 77 372
rect 77 371 78 372
rect 78 371 79 372
rect 79 371 80 372
rect 80 371 81 372
rect 81 371 82 372
rect 82 371 83 372
rect 83 371 84 372
rect 84 371 85 372
rect 85 371 86 372
rect 86 371 87 372
rect 87 371 88 372
rect 88 371 89 372
rect 89 371 90 372
rect 90 371 91 372
rect 148 371 149 372
rect 149 371 150 372
rect 150 371 151 372
rect 151 371 152 372
rect 152 371 153 372
rect 153 371 154 372
rect 154 371 155 372
rect 155 371 156 372
rect 156 371 157 372
rect 157 371 158 372
rect 158 371 159 372
rect 159 371 160 372
rect 160 371 161 372
rect 161 371 162 372
rect 162 371 163 372
rect 163 371 164 372
rect 164 371 165 372
rect 165 371 166 372
rect 334 371 335 372
rect 335 371 336 372
rect 336 371 337 372
rect 337 371 338 372
rect 338 371 339 372
rect 339 371 340 372
rect 340 371 341 372
rect 341 371 342 372
rect 342 371 343 372
rect 343 371 344 372
rect 344 371 345 372
rect 345 371 346 372
rect 346 371 347 372
rect 347 371 348 372
rect 348 371 349 372
rect 349 371 350 372
rect 350 371 351 372
rect 351 371 352 372
rect 352 371 353 372
rect 353 371 354 372
rect 354 371 355 372
rect 355 371 356 372
rect 356 371 357 372
rect 357 371 358 372
rect 358 371 359 372
rect 359 371 360 372
rect 360 371 361 372
rect 361 371 362 372
rect 362 371 363 372
rect 363 371 364 372
rect 364 371 365 372
rect 491 371 492 372
rect 492 371 493 372
rect 493 371 494 372
rect 494 371 495 372
rect 495 371 496 372
rect 496 371 497 372
rect 497 371 498 372
rect 498 371 499 372
rect 499 371 500 372
rect 500 371 501 372
rect 501 371 502 372
rect 502 371 503 372
rect 503 371 504 372
rect 504 371 505 372
rect 505 371 506 372
rect 506 371 507 372
rect 507 371 508 372
rect 508 371 509 372
rect 509 371 510 372
rect 510 371 511 372
rect 511 371 512 372
rect 512 371 513 372
rect 513 371 514 372
rect 514 371 515 372
rect 515 371 516 372
rect 516 371 517 372
rect 517 371 518 372
rect 518 371 519 372
rect 519 371 520 372
rect 520 371 521 372
rect 521 371 522 372
rect 68 370 69 371
rect 69 370 70 371
rect 70 370 71 371
rect 71 370 72 371
rect 72 370 73 371
rect 73 370 74 371
rect 74 370 75 371
rect 75 370 76 371
rect 76 370 77 371
rect 77 370 78 371
rect 78 370 79 371
rect 79 370 80 371
rect 80 370 81 371
rect 81 370 82 371
rect 82 370 83 371
rect 83 370 84 371
rect 84 370 85 371
rect 85 370 86 371
rect 86 370 87 371
rect 87 370 88 371
rect 88 370 89 371
rect 89 370 90 371
rect 90 370 91 371
rect 147 370 148 371
rect 148 370 149 371
rect 149 370 150 371
rect 150 370 151 371
rect 151 370 152 371
rect 152 370 153 371
rect 153 370 154 371
rect 154 370 155 371
rect 155 370 156 371
rect 156 370 157 371
rect 157 370 158 371
rect 158 370 159 371
rect 159 370 160 371
rect 160 370 161 371
rect 161 370 162 371
rect 162 370 163 371
rect 163 370 164 371
rect 164 370 165 371
rect 165 370 166 371
rect 334 370 335 371
rect 335 370 336 371
rect 336 370 337 371
rect 337 370 338 371
rect 338 370 339 371
rect 339 370 340 371
rect 340 370 341 371
rect 341 370 342 371
rect 342 370 343 371
rect 343 370 344 371
rect 344 370 345 371
rect 345 370 346 371
rect 346 370 347 371
rect 347 370 348 371
rect 348 370 349 371
rect 349 370 350 371
rect 350 370 351 371
rect 351 370 352 371
rect 352 370 353 371
rect 353 370 354 371
rect 354 370 355 371
rect 355 370 356 371
rect 356 370 357 371
rect 357 370 358 371
rect 358 370 359 371
rect 359 370 360 371
rect 360 370 361 371
rect 361 370 362 371
rect 362 370 363 371
rect 363 370 364 371
rect 364 370 365 371
rect 491 370 492 371
rect 492 370 493 371
rect 493 370 494 371
rect 494 370 495 371
rect 495 370 496 371
rect 496 370 497 371
rect 497 370 498 371
rect 498 370 499 371
rect 499 370 500 371
rect 500 370 501 371
rect 501 370 502 371
rect 502 370 503 371
rect 503 370 504 371
rect 504 370 505 371
rect 505 370 506 371
rect 506 370 507 371
rect 507 370 508 371
rect 508 370 509 371
rect 509 370 510 371
rect 510 370 511 371
rect 511 370 512 371
rect 512 370 513 371
rect 513 370 514 371
rect 514 370 515 371
rect 515 370 516 371
rect 516 370 517 371
rect 517 370 518 371
rect 518 370 519 371
rect 519 370 520 371
rect 520 370 521 371
rect 521 370 522 371
rect 68 369 69 370
rect 69 369 70 370
rect 70 369 71 370
rect 71 369 72 370
rect 72 369 73 370
rect 73 369 74 370
rect 74 369 75 370
rect 75 369 76 370
rect 76 369 77 370
rect 77 369 78 370
rect 78 369 79 370
rect 79 369 80 370
rect 80 369 81 370
rect 81 369 82 370
rect 82 369 83 370
rect 83 369 84 370
rect 84 369 85 370
rect 85 369 86 370
rect 86 369 87 370
rect 87 369 88 370
rect 147 369 148 370
rect 148 369 149 370
rect 149 369 150 370
rect 150 369 151 370
rect 151 369 152 370
rect 152 369 153 370
rect 153 369 154 370
rect 154 369 155 370
rect 155 369 156 370
rect 156 369 157 370
rect 157 369 158 370
rect 158 369 159 370
rect 159 369 160 370
rect 160 369 161 370
rect 161 369 162 370
rect 162 369 163 370
rect 163 369 164 370
rect 334 369 335 370
rect 335 369 336 370
rect 336 369 337 370
rect 337 369 338 370
rect 338 369 339 370
rect 339 369 340 370
rect 340 369 341 370
rect 341 369 342 370
rect 342 369 343 370
rect 343 369 344 370
rect 344 369 345 370
rect 345 369 346 370
rect 346 369 347 370
rect 347 369 348 370
rect 348 369 349 370
rect 349 369 350 370
rect 350 369 351 370
rect 351 369 352 370
rect 352 369 353 370
rect 353 369 354 370
rect 354 369 355 370
rect 355 369 356 370
rect 356 369 357 370
rect 493 369 494 370
rect 494 369 495 370
rect 495 369 496 370
rect 496 369 497 370
rect 497 369 498 370
rect 498 369 499 370
rect 499 369 500 370
rect 500 369 501 370
rect 501 369 502 370
rect 502 369 503 370
rect 503 369 504 370
rect 504 369 505 370
rect 505 369 506 370
rect 506 369 507 370
rect 507 369 508 370
rect 508 369 509 370
rect 509 369 510 370
rect 510 369 511 370
rect 511 369 512 370
rect 512 369 513 370
rect 513 369 514 370
rect 514 369 515 370
rect 515 369 516 370
rect 516 369 517 370
rect 517 369 518 370
rect 518 369 519 370
rect 519 369 520 370
rect 520 369 521 370
rect 521 369 522 370
rect 66 368 67 369
rect 67 368 68 369
rect 68 368 69 369
rect 69 368 70 369
rect 70 368 71 369
rect 71 368 72 369
rect 72 368 73 369
rect 73 368 74 369
rect 74 368 75 369
rect 75 368 76 369
rect 76 368 77 369
rect 77 368 78 369
rect 78 368 79 369
rect 79 368 80 369
rect 80 368 81 369
rect 81 368 82 369
rect 82 368 83 369
rect 83 368 84 369
rect 84 368 85 369
rect 85 368 86 369
rect 86 368 87 369
rect 87 368 88 369
rect 145 368 146 369
rect 146 368 147 369
rect 147 368 148 369
rect 148 368 149 369
rect 149 368 150 369
rect 150 368 151 369
rect 151 368 152 369
rect 152 368 153 369
rect 153 368 154 369
rect 154 368 155 369
rect 155 368 156 369
rect 156 368 157 369
rect 157 368 158 369
rect 158 368 159 369
rect 159 368 160 369
rect 160 368 161 369
rect 161 368 162 369
rect 162 368 163 369
rect 163 368 164 369
rect 332 368 333 369
rect 333 368 334 369
rect 334 368 335 369
rect 335 368 336 369
rect 336 368 337 369
rect 337 368 338 369
rect 338 368 339 369
rect 339 368 340 369
rect 340 368 341 369
rect 341 368 342 369
rect 342 368 343 369
rect 343 368 344 369
rect 344 368 345 369
rect 345 368 346 369
rect 346 368 347 369
rect 347 368 348 369
rect 348 368 349 369
rect 349 368 350 369
rect 350 368 351 369
rect 351 368 352 369
rect 352 368 353 369
rect 353 368 354 369
rect 354 368 355 369
rect 355 368 356 369
rect 356 368 357 369
rect 493 368 494 369
rect 494 368 495 369
rect 495 368 496 369
rect 496 368 497 369
rect 497 368 498 369
rect 498 368 499 369
rect 499 368 500 369
rect 500 368 501 369
rect 501 368 502 369
rect 502 368 503 369
rect 503 368 504 369
rect 504 368 505 369
rect 505 368 506 369
rect 506 368 507 369
rect 507 368 508 369
rect 508 368 509 369
rect 509 368 510 369
rect 510 368 511 369
rect 511 368 512 369
rect 512 368 513 369
rect 513 368 514 369
rect 514 368 515 369
rect 515 368 516 369
rect 516 368 517 369
rect 517 368 518 369
rect 518 368 519 369
rect 519 368 520 369
rect 520 368 521 369
rect 521 368 522 369
rect 522 368 523 369
rect 523 368 524 369
rect 66 367 67 368
rect 67 367 68 368
rect 68 367 69 368
rect 69 367 70 368
rect 70 367 71 368
rect 71 367 72 368
rect 72 367 73 368
rect 73 367 74 368
rect 74 367 75 368
rect 75 367 76 368
rect 76 367 77 368
rect 77 367 78 368
rect 78 367 79 368
rect 79 367 80 368
rect 80 367 81 368
rect 81 367 82 368
rect 82 367 83 368
rect 83 367 84 368
rect 84 367 85 368
rect 85 367 86 368
rect 145 367 146 368
rect 146 367 147 368
rect 147 367 148 368
rect 148 367 149 368
rect 149 367 150 368
rect 150 367 151 368
rect 151 367 152 368
rect 152 367 153 368
rect 153 367 154 368
rect 154 367 155 368
rect 155 367 156 368
rect 156 367 157 368
rect 157 367 158 368
rect 158 367 159 368
rect 159 367 160 368
rect 160 367 161 368
rect 332 367 333 368
rect 333 367 334 368
rect 334 367 335 368
rect 335 367 336 368
rect 336 367 337 368
rect 337 367 338 368
rect 338 367 339 368
rect 339 367 340 368
rect 340 367 341 368
rect 341 367 342 368
rect 342 367 343 368
rect 343 367 344 368
rect 344 367 345 368
rect 345 367 346 368
rect 346 367 347 368
rect 347 367 348 368
rect 495 367 496 368
rect 496 367 497 368
rect 497 367 498 368
rect 498 367 499 368
rect 499 367 500 368
rect 500 367 501 368
rect 501 367 502 368
rect 502 367 503 368
rect 503 367 504 368
rect 504 367 505 368
rect 505 367 506 368
rect 506 367 507 368
rect 507 367 508 368
rect 508 367 509 368
rect 509 367 510 368
rect 510 367 511 368
rect 511 367 512 368
rect 512 367 513 368
rect 513 367 514 368
rect 514 367 515 368
rect 515 367 516 368
rect 516 367 517 368
rect 517 367 518 368
rect 518 367 519 368
rect 519 367 520 368
rect 520 367 521 368
rect 521 367 522 368
rect 522 367 523 368
rect 523 367 524 368
rect 60 366 61 367
rect 61 366 62 367
rect 62 366 63 367
rect 63 366 64 367
rect 64 366 65 367
rect 65 366 66 367
rect 66 366 67 367
rect 67 366 68 367
rect 68 366 69 367
rect 69 366 70 367
rect 70 366 71 367
rect 71 366 72 367
rect 72 366 73 367
rect 73 366 74 367
rect 74 366 75 367
rect 75 366 76 367
rect 76 366 77 367
rect 77 366 78 367
rect 78 366 79 367
rect 79 366 80 367
rect 80 366 81 367
rect 81 366 82 367
rect 82 366 83 367
rect 83 366 84 367
rect 84 366 85 367
rect 85 366 86 367
rect 143 366 144 367
rect 144 366 145 367
rect 145 366 146 367
rect 146 366 147 367
rect 147 366 148 367
rect 148 366 149 367
rect 149 366 150 367
rect 150 366 151 367
rect 151 366 152 367
rect 152 366 153 367
rect 153 366 154 367
rect 154 366 155 367
rect 155 366 156 367
rect 156 366 157 367
rect 157 366 158 367
rect 158 366 159 367
rect 159 366 160 367
rect 160 366 161 367
rect 330 366 331 367
rect 331 366 332 367
rect 332 366 333 367
rect 333 366 334 367
rect 334 366 335 367
rect 335 366 336 367
rect 336 366 337 367
rect 337 366 338 367
rect 338 366 339 367
rect 339 366 340 367
rect 340 366 341 367
rect 341 366 342 367
rect 342 366 343 367
rect 343 366 344 367
rect 344 366 345 367
rect 345 366 346 367
rect 346 366 347 367
rect 347 366 348 367
rect 495 366 496 367
rect 496 366 497 367
rect 497 366 498 367
rect 498 366 499 367
rect 499 366 500 367
rect 500 366 501 367
rect 501 366 502 367
rect 502 366 503 367
rect 503 366 504 367
rect 504 366 505 367
rect 505 366 506 367
rect 506 366 507 367
rect 507 366 508 367
rect 508 366 509 367
rect 509 366 510 367
rect 510 366 511 367
rect 511 366 512 367
rect 512 366 513 367
rect 513 366 514 367
rect 514 366 515 367
rect 515 366 516 367
rect 516 366 517 367
rect 517 366 518 367
rect 518 366 519 367
rect 519 366 520 367
rect 520 366 521 367
rect 521 366 522 367
rect 522 366 523 367
rect 523 366 524 367
rect 524 366 525 367
rect 525 366 526 367
rect 60 365 61 366
rect 61 365 62 366
rect 62 365 63 366
rect 63 365 64 366
rect 64 365 65 366
rect 65 365 66 366
rect 66 365 67 366
rect 67 365 68 366
rect 68 365 69 366
rect 69 365 70 366
rect 70 365 71 366
rect 71 365 72 366
rect 72 365 73 366
rect 73 365 74 366
rect 74 365 75 366
rect 75 365 76 366
rect 76 365 77 366
rect 77 365 78 366
rect 78 365 79 366
rect 79 365 80 366
rect 143 365 144 366
rect 144 365 145 366
rect 145 365 146 366
rect 146 365 147 366
rect 147 365 148 366
rect 148 365 149 366
rect 149 365 150 366
rect 150 365 151 366
rect 151 365 152 366
rect 152 365 153 366
rect 153 365 154 366
rect 154 365 155 366
rect 155 365 156 366
rect 156 365 157 366
rect 157 365 158 366
rect 158 365 159 366
rect 159 365 160 366
rect 160 365 161 366
rect 330 365 331 366
rect 331 365 332 366
rect 332 365 333 366
rect 336 365 337 366
rect 337 365 338 366
rect 338 365 339 366
rect 497 365 498 366
rect 498 365 499 366
rect 499 365 500 366
rect 500 365 501 366
rect 501 365 502 366
rect 502 365 503 366
rect 503 365 504 366
rect 504 365 505 366
rect 505 365 506 366
rect 506 365 507 366
rect 507 365 508 366
rect 508 365 509 366
rect 509 365 510 366
rect 510 365 511 366
rect 511 365 512 366
rect 512 365 513 366
rect 513 365 514 366
rect 514 365 515 366
rect 515 365 516 366
rect 516 365 517 366
rect 517 365 518 366
rect 518 365 519 366
rect 519 365 520 366
rect 520 365 521 366
rect 521 365 522 366
rect 522 365 523 366
rect 523 365 524 366
rect 524 365 525 366
rect 525 365 526 366
rect 57 364 58 365
rect 58 364 59 365
rect 59 364 60 365
rect 60 364 61 365
rect 61 364 62 365
rect 62 364 63 365
rect 63 364 64 365
rect 64 364 65 365
rect 65 364 66 365
rect 66 364 67 365
rect 67 364 68 365
rect 68 364 69 365
rect 69 364 70 365
rect 70 364 71 365
rect 71 364 72 365
rect 72 364 73 365
rect 73 364 74 365
rect 74 364 75 365
rect 75 364 76 365
rect 76 364 77 365
rect 77 364 78 365
rect 78 364 79 365
rect 79 364 80 365
rect 141 364 142 365
rect 142 364 143 365
rect 143 364 144 365
rect 144 364 145 365
rect 145 364 146 365
rect 146 364 147 365
rect 147 364 148 365
rect 148 364 149 365
rect 149 364 150 365
rect 150 364 151 365
rect 151 364 152 365
rect 152 364 153 365
rect 153 364 154 365
rect 154 364 155 365
rect 155 364 156 365
rect 156 364 157 365
rect 157 364 158 365
rect 158 364 159 365
rect 159 364 160 365
rect 160 364 161 365
rect 330 364 331 365
rect 331 364 332 365
rect 332 364 333 365
rect 336 364 337 365
rect 337 364 338 365
rect 338 364 339 365
rect 497 364 498 365
rect 498 364 499 365
rect 499 364 500 365
rect 500 364 501 365
rect 501 364 502 365
rect 502 364 503 365
rect 503 364 504 365
rect 504 364 505 365
rect 505 364 506 365
rect 506 364 507 365
rect 507 364 508 365
rect 508 364 509 365
rect 509 364 510 365
rect 510 364 511 365
rect 511 364 512 365
rect 512 364 513 365
rect 513 364 514 365
rect 514 364 515 365
rect 515 364 516 365
rect 516 364 517 365
rect 517 364 518 365
rect 518 364 519 365
rect 519 364 520 365
rect 520 364 521 365
rect 521 364 522 365
rect 522 364 523 365
rect 523 364 524 365
rect 524 364 525 365
rect 525 364 526 365
rect 57 363 58 364
rect 58 363 59 364
rect 59 363 60 364
rect 60 363 61 364
rect 61 363 62 364
rect 62 363 63 364
rect 63 363 64 364
rect 64 363 65 364
rect 65 363 66 364
rect 66 363 67 364
rect 67 363 68 364
rect 68 363 69 364
rect 69 363 70 364
rect 70 363 71 364
rect 71 363 72 364
rect 72 363 73 364
rect 73 363 74 364
rect 74 363 75 364
rect 75 363 76 364
rect 141 363 142 364
rect 142 363 143 364
rect 143 363 144 364
rect 144 363 145 364
rect 145 363 146 364
rect 146 363 147 364
rect 147 363 148 364
rect 148 363 149 364
rect 149 363 150 364
rect 150 363 151 364
rect 151 363 152 364
rect 152 363 153 364
rect 153 363 154 364
rect 154 363 155 364
rect 155 363 156 364
rect 156 363 157 364
rect 499 363 500 364
rect 500 363 501 364
rect 501 363 502 364
rect 502 363 503 364
rect 503 363 504 364
rect 504 363 505 364
rect 505 363 506 364
rect 506 363 507 364
rect 507 363 508 364
rect 508 363 509 364
rect 509 363 510 364
rect 510 363 511 364
rect 511 363 512 364
rect 512 363 513 364
rect 513 363 514 364
rect 514 363 515 364
rect 515 363 516 364
rect 516 363 517 364
rect 517 363 518 364
rect 518 363 519 364
rect 519 363 520 364
rect 520 363 521 364
rect 521 363 522 364
rect 522 363 523 364
rect 523 363 524 364
rect 524 363 525 364
rect 525 363 526 364
rect 53 362 54 363
rect 54 362 55 363
rect 55 362 56 363
rect 56 362 57 363
rect 57 362 58 363
rect 58 362 59 363
rect 59 362 60 363
rect 60 362 61 363
rect 61 362 62 363
rect 62 362 63 363
rect 63 362 64 363
rect 64 362 65 363
rect 65 362 66 363
rect 66 362 67 363
rect 67 362 68 363
rect 68 362 69 363
rect 69 362 70 363
rect 70 362 71 363
rect 71 362 72 363
rect 72 362 73 363
rect 73 362 74 363
rect 74 362 75 363
rect 75 362 76 363
rect 139 362 140 363
rect 140 362 141 363
rect 141 362 142 363
rect 142 362 143 363
rect 143 362 144 363
rect 144 362 145 363
rect 145 362 146 363
rect 146 362 147 363
rect 147 362 148 363
rect 148 362 149 363
rect 149 362 150 363
rect 150 362 151 363
rect 151 362 152 363
rect 152 362 153 363
rect 153 362 154 363
rect 154 362 155 363
rect 155 362 156 363
rect 156 362 157 363
rect 499 362 500 363
rect 500 362 501 363
rect 501 362 502 363
rect 502 362 503 363
rect 503 362 504 363
rect 504 362 505 363
rect 505 362 506 363
rect 506 362 507 363
rect 507 362 508 363
rect 508 362 509 363
rect 509 362 510 363
rect 510 362 511 363
rect 511 362 512 363
rect 512 362 513 363
rect 513 362 514 363
rect 514 362 515 363
rect 515 362 516 363
rect 516 362 517 363
rect 517 362 518 363
rect 518 362 519 363
rect 519 362 520 363
rect 520 362 521 363
rect 521 362 522 363
rect 522 362 523 363
rect 523 362 524 363
rect 524 362 525 363
rect 525 362 526 363
rect 526 362 527 363
rect 527 362 528 363
rect 53 361 54 362
rect 54 361 55 362
rect 55 361 56 362
rect 56 361 57 362
rect 57 361 58 362
rect 58 361 59 362
rect 59 361 60 362
rect 60 361 61 362
rect 61 361 62 362
rect 62 361 63 362
rect 63 361 64 362
rect 64 361 65 362
rect 65 361 66 362
rect 66 361 67 362
rect 67 361 68 362
rect 68 361 69 362
rect 69 361 70 362
rect 70 361 71 362
rect 71 361 72 362
rect 72 361 73 362
rect 73 361 74 362
rect 139 361 140 362
rect 140 361 141 362
rect 141 361 142 362
rect 142 361 143 362
rect 143 361 144 362
rect 144 361 145 362
rect 145 361 146 362
rect 146 361 147 362
rect 147 361 148 362
rect 148 361 149 362
rect 149 361 150 362
rect 150 361 151 362
rect 151 361 152 362
rect 152 361 153 362
rect 153 361 154 362
rect 154 361 155 362
rect 155 361 156 362
rect 156 361 157 362
rect 499 361 500 362
rect 500 361 501 362
rect 501 361 502 362
rect 502 361 503 362
rect 503 361 504 362
rect 504 361 505 362
rect 505 361 506 362
rect 506 361 507 362
rect 507 361 508 362
rect 508 361 509 362
rect 509 361 510 362
rect 510 361 511 362
rect 511 361 512 362
rect 512 361 513 362
rect 513 361 514 362
rect 514 361 515 362
rect 515 361 516 362
rect 516 361 517 362
rect 517 361 518 362
rect 518 361 519 362
rect 519 361 520 362
rect 520 361 521 362
rect 521 361 522 362
rect 522 361 523 362
rect 523 361 524 362
rect 524 361 525 362
rect 525 361 526 362
rect 526 361 527 362
rect 527 361 528 362
rect 47 360 48 361
rect 48 360 49 361
rect 49 360 50 361
rect 50 360 51 361
rect 51 360 52 361
rect 52 360 53 361
rect 53 360 54 361
rect 54 360 55 361
rect 55 360 56 361
rect 56 360 57 361
rect 57 360 58 361
rect 58 360 59 361
rect 59 360 60 361
rect 60 360 61 361
rect 61 360 62 361
rect 62 360 63 361
rect 63 360 64 361
rect 64 360 65 361
rect 65 360 66 361
rect 66 360 67 361
rect 67 360 68 361
rect 68 360 69 361
rect 69 360 70 361
rect 70 360 71 361
rect 71 360 72 361
rect 72 360 73 361
rect 73 360 74 361
rect 137 360 138 361
rect 138 360 139 361
rect 139 360 140 361
rect 140 360 141 361
rect 141 360 142 361
rect 142 360 143 361
rect 143 360 144 361
rect 144 360 145 361
rect 145 360 146 361
rect 146 360 147 361
rect 147 360 148 361
rect 148 360 149 361
rect 149 360 150 361
rect 150 360 151 361
rect 151 360 152 361
rect 152 360 153 361
rect 153 360 154 361
rect 154 360 155 361
rect 155 360 156 361
rect 156 360 157 361
rect 499 360 500 361
rect 500 360 501 361
rect 501 360 502 361
rect 502 360 503 361
rect 503 360 504 361
rect 504 360 505 361
rect 505 360 506 361
rect 506 360 507 361
rect 507 360 508 361
rect 508 360 509 361
rect 509 360 510 361
rect 510 360 511 361
rect 511 360 512 361
rect 512 360 513 361
rect 513 360 514 361
rect 514 360 515 361
rect 515 360 516 361
rect 516 360 517 361
rect 517 360 518 361
rect 518 360 519 361
rect 519 360 520 361
rect 520 360 521 361
rect 521 360 522 361
rect 522 360 523 361
rect 523 360 524 361
rect 524 360 525 361
rect 525 360 526 361
rect 526 360 527 361
rect 527 360 528 361
rect 47 359 48 360
rect 48 359 49 360
rect 49 359 50 360
rect 50 359 51 360
rect 51 359 52 360
rect 52 359 53 360
rect 53 359 54 360
rect 54 359 55 360
rect 55 359 56 360
rect 56 359 57 360
rect 57 359 58 360
rect 58 359 59 360
rect 59 359 60 360
rect 60 359 61 360
rect 61 359 62 360
rect 62 359 63 360
rect 63 359 64 360
rect 64 359 65 360
rect 65 359 66 360
rect 66 359 67 360
rect 67 359 68 360
rect 68 359 69 360
rect 137 359 138 360
rect 138 359 139 360
rect 139 359 140 360
rect 140 359 141 360
rect 141 359 142 360
rect 142 359 143 360
rect 143 359 144 360
rect 144 359 145 360
rect 145 359 146 360
rect 146 359 147 360
rect 147 359 148 360
rect 148 359 149 360
rect 149 359 150 360
rect 150 359 151 360
rect 151 359 152 360
rect 152 359 153 360
rect 153 359 154 360
rect 154 359 155 360
rect 501 359 502 360
rect 502 359 503 360
rect 503 359 504 360
rect 504 359 505 360
rect 505 359 506 360
rect 506 359 507 360
rect 507 359 508 360
rect 508 359 509 360
rect 509 359 510 360
rect 510 359 511 360
rect 511 359 512 360
rect 512 359 513 360
rect 513 359 514 360
rect 514 359 515 360
rect 515 359 516 360
rect 516 359 517 360
rect 517 359 518 360
rect 518 359 519 360
rect 519 359 520 360
rect 520 359 521 360
rect 521 359 522 360
rect 522 359 523 360
rect 523 359 524 360
rect 524 359 525 360
rect 525 359 526 360
rect 526 359 527 360
rect 527 359 528 360
rect 44 358 45 359
rect 45 358 46 359
rect 46 358 47 359
rect 47 358 48 359
rect 48 358 49 359
rect 49 358 50 359
rect 50 358 51 359
rect 51 358 52 359
rect 52 358 53 359
rect 53 358 54 359
rect 54 358 55 359
rect 55 358 56 359
rect 56 358 57 359
rect 57 358 58 359
rect 58 358 59 359
rect 59 358 60 359
rect 60 358 61 359
rect 61 358 62 359
rect 62 358 63 359
rect 63 358 64 359
rect 64 358 65 359
rect 65 358 66 359
rect 66 358 67 359
rect 67 358 68 359
rect 68 358 69 359
rect 135 358 136 359
rect 136 358 137 359
rect 137 358 138 359
rect 138 358 139 359
rect 139 358 140 359
rect 140 358 141 359
rect 141 358 142 359
rect 142 358 143 359
rect 143 358 144 359
rect 144 358 145 359
rect 145 358 146 359
rect 146 358 147 359
rect 147 358 148 359
rect 148 358 149 359
rect 149 358 150 359
rect 150 358 151 359
rect 151 358 152 359
rect 152 358 153 359
rect 153 358 154 359
rect 154 358 155 359
rect 501 358 502 359
rect 502 358 503 359
rect 503 358 504 359
rect 504 358 505 359
rect 505 358 506 359
rect 506 358 507 359
rect 507 358 508 359
rect 508 358 509 359
rect 509 358 510 359
rect 510 358 511 359
rect 511 358 512 359
rect 512 358 513 359
rect 513 358 514 359
rect 514 358 515 359
rect 515 358 516 359
rect 516 358 517 359
rect 517 358 518 359
rect 518 358 519 359
rect 519 358 520 359
rect 520 358 521 359
rect 521 358 522 359
rect 522 358 523 359
rect 523 358 524 359
rect 524 358 525 359
rect 525 358 526 359
rect 526 358 527 359
rect 527 358 528 359
rect 528 358 529 359
rect 529 358 530 359
rect 44 357 45 358
rect 45 357 46 358
rect 46 357 47 358
rect 47 357 48 358
rect 48 357 49 358
rect 49 357 50 358
rect 50 357 51 358
rect 51 357 52 358
rect 52 357 53 358
rect 53 357 54 358
rect 54 357 55 358
rect 55 357 56 358
rect 56 357 57 358
rect 57 357 58 358
rect 58 357 59 358
rect 59 357 60 358
rect 60 357 61 358
rect 61 357 62 358
rect 62 357 63 358
rect 135 357 136 358
rect 136 357 137 358
rect 137 357 138 358
rect 138 357 139 358
rect 139 357 140 358
rect 140 357 141 358
rect 141 357 142 358
rect 142 357 143 358
rect 143 357 144 358
rect 144 357 145 358
rect 145 357 146 358
rect 146 357 147 358
rect 147 357 148 358
rect 148 357 149 358
rect 149 357 150 358
rect 150 357 151 358
rect 502 357 503 358
rect 503 357 504 358
rect 504 357 505 358
rect 505 357 506 358
rect 506 357 507 358
rect 507 357 508 358
rect 508 357 509 358
rect 509 357 510 358
rect 510 357 511 358
rect 511 357 512 358
rect 512 357 513 358
rect 513 357 514 358
rect 514 357 515 358
rect 515 357 516 358
rect 516 357 517 358
rect 517 357 518 358
rect 518 357 519 358
rect 519 357 520 358
rect 520 357 521 358
rect 521 357 522 358
rect 522 357 523 358
rect 523 357 524 358
rect 524 357 525 358
rect 525 357 526 358
rect 526 357 527 358
rect 527 357 528 358
rect 528 357 529 358
rect 529 357 530 358
rect 40 356 41 357
rect 41 356 42 357
rect 42 356 43 357
rect 43 356 44 357
rect 44 356 45 357
rect 45 356 46 357
rect 46 356 47 357
rect 47 356 48 357
rect 48 356 49 357
rect 49 356 50 357
rect 50 356 51 357
rect 51 356 52 357
rect 52 356 53 357
rect 53 356 54 357
rect 54 356 55 357
rect 55 356 56 357
rect 56 356 57 357
rect 57 356 58 357
rect 58 356 59 357
rect 59 356 60 357
rect 60 356 61 357
rect 61 356 62 357
rect 62 356 63 357
rect 133 356 134 357
rect 134 356 135 357
rect 135 356 136 357
rect 136 356 137 357
rect 137 356 138 357
rect 138 356 139 357
rect 139 356 140 357
rect 140 356 141 357
rect 141 356 142 357
rect 142 356 143 357
rect 143 356 144 357
rect 144 356 145 357
rect 145 356 146 357
rect 146 356 147 357
rect 147 356 148 357
rect 148 356 149 357
rect 149 356 150 357
rect 150 356 151 357
rect 502 356 503 357
rect 503 356 504 357
rect 504 356 505 357
rect 505 356 506 357
rect 506 356 507 357
rect 507 356 508 357
rect 508 356 509 357
rect 509 356 510 357
rect 510 356 511 357
rect 511 356 512 357
rect 512 356 513 357
rect 513 356 514 357
rect 514 356 515 357
rect 515 356 516 357
rect 516 356 517 357
rect 517 356 518 357
rect 518 356 519 357
rect 519 356 520 357
rect 520 356 521 357
rect 521 356 522 357
rect 522 356 523 357
rect 523 356 524 357
rect 524 356 525 357
rect 525 356 526 357
rect 526 356 527 357
rect 527 356 528 357
rect 528 356 529 357
rect 529 356 530 357
rect 40 355 41 356
rect 41 355 42 356
rect 42 355 43 356
rect 43 355 44 356
rect 44 355 45 356
rect 45 355 46 356
rect 46 355 47 356
rect 47 355 48 356
rect 48 355 49 356
rect 49 355 50 356
rect 50 355 51 356
rect 51 355 52 356
rect 52 355 53 356
rect 53 355 54 356
rect 54 355 55 356
rect 55 355 56 356
rect 56 355 57 356
rect 57 355 58 356
rect 58 355 59 356
rect 133 355 134 356
rect 134 355 135 356
rect 135 355 136 356
rect 136 355 137 356
rect 137 355 138 356
rect 138 355 139 356
rect 139 355 140 356
rect 140 355 141 356
rect 141 355 142 356
rect 142 355 143 356
rect 143 355 144 356
rect 144 355 145 356
rect 145 355 146 356
rect 146 355 147 356
rect 147 355 148 356
rect 148 355 149 356
rect 149 355 150 356
rect 150 355 151 356
rect 504 355 505 356
rect 505 355 506 356
rect 506 355 507 356
rect 507 355 508 356
rect 508 355 509 356
rect 509 355 510 356
rect 510 355 511 356
rect 511 355 512 356
rect 512 355 513 356
rect 513 355 514 356
rect 514 355 515 356
rect 515 355 516 356
rect 516 355 517 356
rect 517 355 518 356
rect 518 355 519 356
rect 519 355 520 356
rect 520 355 521 356
rect 521 355 522 356
rect 522 355 523 356
rect 523 355 524 356
rect 524 355 525 356
rect 525 355 526 356
rect 526 355 527 356
rect 527 355 528 356
rect 528 355 529 356
rect 529 355 530 356
rect 36 354 37 355
rect 37 354 38 355
rect 38 354 39 355
rect 39 354 40 355
rect 40 354 41 355
rect 41 354 42 355
rect 42 354 43 355
rect 43 354 44 355
rect 44 354 45 355
rect 45 354 46 355
rect 46 354 47 355
rect 47 354 48 355
rect 48 354 49 355
rect 49 354 50 355
rect 50 354 51 355
rect 51 354 52 355
rect 52 354 53 355
rect 53 354 54 355
rect 54 354 55 355
rect 55 354 56 355
rect 56 354 57 355
rect 57 354 58 355
rect 58 354 59 355
rect 132 354 133 355
rect 133 354 134 355
rect 134 354 135 355
rect 135 354 136 355
rect 136 354 137 355
rect 137 354 138 355
rect 138 354 139 355
rect 139 354 140 355
rect 140 354 141 355
rect 141 354 142 355
rect 142 354 143 355
rect 143 354 144 355
rect 144 354 145 355
rect 145 354 146 355
rect 146 354 147 355
rect 147 354 148 355
rect 148 354 149 355
rect 149 354 150 355
rect 150 354 151 355
rect 504 354 505 355
rect 505 354 506 355
rect 506 354 507 355
rect 507 354 508 355
rect 508 354 509 355
rect 509 354 510 355
rect 510 354 511 355
rect 511 354 512 355
rect 512 354 513 355
rect 513 354 514 355
rect 514 354 515 355
rect 515 354 516 355
rect 516 354 517 355
rect 517 354 518 355
rect 518 354 519 355
rect 519 354 520 355
rect 520 354 521 355
rect 521 354 522 355
rect 522 354 523 355
rect 523 354 524 355
rect 524 354 525 355
rect 525 354 526 355
rect 526 354 527 355
rect 527 354 528 355
rect 528 354 529 355
rect 529 354 530 355
rect 36 353 37 354
rect 37 353 38 354
rect 38 353 39 354
rect 39 353 40 354
rect 40 353 41 354
rect 41 353 42 354
rect 42 353 43 354
rect 43 353 44 354
rect 44 353 45 354
rect 45 353 46 354
rect 46 353 47 354
rect 47 353 48 354
rect 48 353 49 354
rect 49 353 50 354
rect 50 353 51 354
rect 51 353 52 354
rect 52 353 53 354
rect 53 353 54 354
rect 132 353 133 354
rect 133 353 134 354
rect 134 353 135 354
rect 135 353 136 354
rect 136 353 137 354
rect 137 353 138 354
rect 138 353 139 354
rect 139 353 140 354
rect 140 353 141 354
rect 141 353 142 354
rect 142 353 143 354
rect 143 353 144 354
rect 144 353 145 354
rect 145 353 146 354
rect 146 353 147 354
rect 147 353 148 354
rect 148 353 149 354
rect 504 353 505 354
rect 505 353 506 354
rect 506 353 507 354
rect 507 353 508 354
rect 508 353 509 354
rect 509 353 510 354
rect 510 353 511 354
rect 511 353 512 354
rect 512 353 513 354
rect 513 353 514 354
rect 514 353 515 354
rect 515 353 516 354
rect 516 353 517 354
rect 517 353 518 354
rect 518 353 519 354
rect 519 353 520 354
rect 520 353 521 354
rect 521 353 522 354
rect 522 353 523 354
rect 523 353 524 354
rect 524 353 525 354
rect 525 353 526 354
rect 526 353 527 354
rect 527 353 528 354
rect 528 353 529 354
rect 529 353 530 354
rect 30 352 31 353
rect 31 352 32 353
rect 32 352 33 353
rect 33 352 34 353
rect 34 352 35 353
rect 35 352 36 353
rect 36 352 37 353
rect 37 352 38 353
rect 38 352 39 353
rect 39 352 40 353
rect 40 352 41 353
rect 41 352 42 353
rect 42 352 43 353
rect 43 352 44 353
rect 44 352 45 353
rect 45 352 46 353
rect 46 352 47 353
rect 47 352 48 353
rect 48 352 49 353
rect 49 352 50 353
rect 50 352 51 353
rect 51 352 52 353
rect 52 352 53 353
rect 53 352 54 353
rect 130 352 131 353
rect 131 352 132 353
rect 132 352 133 353
rect 133 352 134 353
rect 134 352 135 353
rect 135 352 136 353
rect 136 352 137 353
rect 137 352 138 353
rect 138 352 139 353
rect 139 352 140 353
rect 140 352 141 353
rect 141 352 142 353
rect 142 352 143 353
rect 143 352 144 353
rect 144 352 145 353
rect 145 352 146 353
rect 146 352 147 353
rect 147 352 148 353
rect 148 352 149 353
rect 504 352 505 353
rect 505 352 506 353
rect 506 352 507 353
rect 507 352 508 353
rect 508 352 509 353
rect 509 352 510 353
rect 510 352 511 353
rect 511 352 512 353
rect 512 352 513 353
rect 513 352 514 353
rect 514 352 515 353
rect 515 352 516 353
rect 516 352 517 353
rect 517 352 518 353
rect 518 352 519 353
rect 519 352 520 353
rect 520 352 521 353
rect 521 352 522 353
rect 522 352 523 353
rect 523 352 524 353
rect 524 352 525 353
rect 525 352 526 353
rect 526 352 527 353
rect 527 352 528 353
rect 528 352 529 353
rect 529 352 530 353
rect 530 352 531 353
rect 30 351 31 352
rect 31 351 32 352
rect 32 351 33 352
rect 33 351 34 352
rect 34 351 35 352
rect 35 351 36 352
rect 36 351 37 352
rect 37 351 38 352
rect 38 351 39 352
rect 39 351 40 352
rect 40 351 41 352
rect 41 351 42 352
rect 42 351 43 352
rect 43 351 44 352
rect 44 351 45 352
rect 45 351 46 352
rect 130 351 131 352
rect 131 351 132 352
rect 132 351 133 352
rect 133 351 134 352
rect 134 351 135 352
rect 135 351 136 352
rect 136 351 137 352
rect 137 351 138 352
rect 138 351 139 352
rect 139 351 140 352
rect 140 351 141 352
rect 141 351 142 352
rect 142 351 143 352
rect 143 351 144 352
rect 144 351 145 352
rect 145 351 146 352
rect 506 351 507 352
rect 507 351 508 352
rect 508 351 509 352
rect 509 351 510 352
rect 510 351 511 352
rect 511 351 512 352
rect 512 351 513 352
rect 513 351 514 352
rect 514 351 515 352
rect 515 351 516 352
rect 516 351 517 352
rect 517 351 518 352
rect 518 351 519 352
rect 519 351 520 352
rect 520 351 521 352
rect 521 351 522 352
rect 522 351 523 352
rect 523 351 524 352
rect 524 351 525 352
rect 525 351 526 352
rect 526 351 527 352
rect 527 351 528 352
rect 528 351 529 352
rect 529 351 530 352
rect 530 351 531 352
rect 27 350 28 351
rect 28 350 29 351
rect 29 350 30 351
rect 30 350 31 351
rect 31 350 32 351
rect 32 350 33 351
rect 33 350 34 351
rect 34 350 35 351
rect 35 350 36 351
rect 36 350 37 351
rect 37 350 38 351
rect 38 350 39 351
rect 39 350 40 351
rect 40 350 41 351
rect 41 350 42 351
rect 42 350 43 351
rect 43 350 44 351
rect 44 350 45 351
rect 45 350 46 351
rect 128 350 129 351
rect 129 350 130 351
rect 130 350 131 351
rect 131 350 132 351
rect 132 350 133 351
rect 133 350 134 351
rect 134 350 135 351
rect 135 350 136 351
rect 136 350 137 351
rect 137 350 138 351
rect 138 350 139 351
rect 139 350 140 351
rect 140 350 141 351
rect 141 350 142 351
rect 142 350 143 351
rect 143 350 144 351
rect 144 350 145 351
rect 145 350 146 351
rect 506 350 507 351
rect 507 350 508 351
rect 508 350 509 351
rect 509 350 510 351
rect 510 350 511 351
rect 511 350 512 351
rect 512 350 513 351
rect 513 350 514 351
rect 514 350 515 351
rect 515 350 516 351
rect 516 350 517 351
rect 517 350 518 351
rect 518 350 519 351
rect 519 350 520 351
rect 520 350 521 351
rect 521 350 522 351
rect 522 350 523 351
rect 523 350 524 351
rect 524 350 525 351
rect 525 350 526 351
rect 526 350 527 351
rect 527 350 528 351
rect 528 350 529 351
rect 529 350 530 351
rect 530 350 531 351
rect 27 349 28 350
rect 28 349 29 350
rect 29 349 30 350
rect 30 349 31 350
rect 31 349 32 350
rect 32 349 33 350
rect 33 349 34 350
rect 34 349 35 350
rect 35 349 36 350
rect 36 349 37 350
rect 37 349 38 350
rect 38 349 39 350
rect 39 349 40 350
rect 40 349 41 350
rect 41 349 42 350
rect 42 349 43 350
rect 128 349 129 350
rect 129 349 130 350
rect 130 349 131 350
rect 131 349 132 350
rect 132 349 133 350
rect 133 349 134 350
rect 134 349 135 350
rect 135 349 136 350
rect 136 349 137 350
rect 137 349 138 350
rect 138 349 139 350
rect 139 349 140 350
rect 140 349 141 350
rect 141 349 142 350
rect 142 349 143 350
rect 143 349 144 350
rect 144 349 145 350
rect 145 349 146 350
rect 508 349 509 350
rect 509 349 510 350
rect 510 349 511 350
rect 511 349 512 350
rect 512 349 513 350
rect 513 349 514 350
rect 514 349 515 350
rect 515 349 516 350
rect 516 349 517 350
rect 517 349 518 350
rect 518 349 519 350
rect 519 349 520 350
rect 520 349 521 350
rect 521 349 522 350
rect 522 349 523 350
rect 523 349 524 350
rect 524 349 525 350
rect 525 349 526 350
rect 526 349 527 350
rect 527 349 528 350
rect 528 349 529 350
rect 529 349 530 350
rect 530 349 531 350
rect 23 348 24 349
rect 24 348 25 349
rect 25 348 26 349
rect 26 348 27 349
rect 27 348 28 349
rect 28 348 29 349
rect 29 348 30 349
rect 30 348 31 349
rect 31 348 32 349
rect 32 348 33 349
rect 33 348 34 349
rect 34 348 35 349
rect 35 348 36 349
rect 36 348 37 349
rect 37 348 38 349
rect 38 348 39 349
rect 39 348 40 349
rect 40 348 41 349
rect 41 348 42 349
rect 42 348 43 349
rect 126 348 127 349
rect 127 348 128 349
rect 128 348 129 349
rect 129 348 130 349
rect 130 348 131 349
rect 131 348 132 349
rect 132 348 133 349
rect 133 348 134 349
rect 134 348 135 349
rect 135 348 136 349
rect 136 348 137 349
rect 137 348 138 349
rect 138 348 139 349
rect 139 348 140 349
rect 140 348 141 349
rect 141 348 142 349
rect 142 348 143 349
rect 143 348 144 349
rect 144 348 145 349
rect 145 348 146 349
rect 508 348 509 349
rect 509 348 510 349
rect 510 348 511 349
rect 511 348 512 349
rect 512 348 513 349
rect 513 348 514 349
rect 514 348 515 349
rect 515 348 516 349
rect 516 348 517 349
rect 517 348 518 349
rect 518 348 519 349
rect 519 348 520 349
rect 520 348 521 349
rect 521 348 522 349
rect 522 348 523 349
rect 523 348 524 349
rect 524 348 525 349
rect 525 348 526 349
rect 526 348 527 349
rect 527 348 528 349
rect 528 348 529 349
rect 529 348 530 349
rect 530 348 531 349
rect 23 347 24 348
rect 24 347 25 348
rect 25 347 26 348
rect 26 347 27 348
rect 27 347 28 348
rect 28 347 29 348
rect 29 347 30 348
rect 30 347 31 348
rect 31 347 32 348
rect 32 347 33 348
rect 33 347 34 348
rect 34 347 35 348
rect 126 347 127 348
rect 127 347 128 348
rect 128 347 129 348
rect 129 347 130 348
rect 130 347 131 348
rect 131 347 132 348
rect 132 347 133 348
rect 133 347 134 348
rect 134 347 135 348
rect 135 347 136 348
rect 136 347 137 348
rect 137 347 138 348
rect 138 347 139 348
rect 139 347 140 348
rect 140 347 141 348
rect 141 347 142 348
rect 142 347 143 348
rect 143 347 144 348
rect 508 347 509 348
rect 509 347 510 348
rect 510 347 511 348
rect 511 347 512 348
rect 512 347 513 348
rect 513 347 514 348
rect 514 347 515 348
rect 515 347 516 348
rect 516 347 517 348
rect 517 347 518 348
rect 518 347 519 348
rect 519 347 520 348
rect 520 347 521 348
rect 521 347 522 348
rect 522 347 523 348
rect 523 347 524 348
rect 524 347 525 348
rect 525 347 526 348
rect 526 347 527 348
rect 527 347 528 348
rect 528 347 529 348
rect 529 347 530 348
rect 530 347 531 348
rect 21 346 22 347
rect 22 346 23 347
rect 23 346 24 347
rect 24 346 25 347
rect 25 346 26 347
rect 26 346 27 347
rect 27 346 28 347
rect 28 346 29 347
rect 29 346 30 347
rect 30 346 31 347
rect 31 346 32 347
rect 32 346 33 347
rect 33 346 34 347
rect 34 346 35 347
rect 124 346 125 347
rect 125 346 126 347
rect 126 346 127 347
rect 127 346 128 347
rect 128 346 129 347
rect 129 346 130 347
rect 130 346 131 347
rect 131 346 132 347
rect 132 346 133 347
rect 133 346 134 347
rect 134 346 135 347
rect 135 346 136 347
rect 136 346 137 347
rect 137 346 138 347
rect 138 346 139 347
rect 139 346 140 347
rect 140 346 141 347
rect 141 346 142 347
rect 142 346 143 347
rect 143 346 144 347
rect 508 346 509 347
rect 509 346 510 347
rect 510 346 511 347
rect 511 346 512 347
rect 512 346 513 347
rect 513 346 514 347
rect 514 346 515 347
rect 515 346 516 347
rect 516 346 517 347
rect 517 346 518 347
rect 518 346 519 347
rect 519 346 520 347
rect 520 346 521 347
rect 521 346 522 347
rect 522 346 523 347
rect 523 346 524 347
rect 524 346 525 347
rect 525 346 526 347
rect 526 346 527 347
rect 527 346 528 347
rect 528 346 529 347
rect 529 346 530 347
rect 530 346 531 347
rect 531 346 532 347
rect 532 346 533 347
rect 21 345 22 346
rect 22 345 23 346
rect 23 345 24 346
rect 24 345 25 346
rect 25 345 26 346
rect 26 345 27 346
rect 27 345 28 346
rect 28 345 29 346
rect 29 345 30 346
rect 124 345 125 346
rect 125 345 126 346
rect 126 345 127 346
rect 127 345 128 346
rect 128 345 129 346
rect 129 345 130 346
rect 130 345 131 346
rect 131 345 132 346
rect 132 345 133 346
rect 133 345 134 346
rect 134 345 135 346
rect 135 345 136 346
rect 136 345 137 346
rect 137 345 138 346
rect 138 345 139 346
rect 139 345 140 346
rect 510 345 511 346
rect 511 345 512 346
rect 512 345 513 346
rect 513 345 514 346
rect 514 345 515 346
rect 515 345 516 346
rect 516 345 517 346
rect 517 345 518 346
rect 518 345 519 346
rect 519 345 520 346
rect 520 345 521 346
rect 521 345 522 346
rect 522 345 523 346
rect 523 345 524 346
rect 524 345 525 346
rect 525 345 526 346
rect 526 345 527 346
rect 527 345 528 346
rect 528 345 529 346
rect 529 345 530 346
rect 530 345 531 346
rect 531 345 532 346
rect 532 345 533 346
rect 21 344 22 345
rect 22 344 23 345
rect 23 344 24 345
rect 24 344 25 345
rect 25 344 26 345
rect 26 344 27 345
rect 27 344 28 345
rect 28 344 29 345
rect 29 344 30 345
rect 30 344 31 345
rect 122 344 123 345
rect 123 344 124 345
rect 124 344 125 345
rect 125 344 126 345
rect 126 344 127 345
rect 127 344 128 345
rect 128 344 129 345
rect 129 344 130 345
rect 130 344 131 345
rect 131 344 132 345
rect 132 344 133 345
rect 133 344 134 345
rect 134 344 135 345
rect 135 344 136 345
rect 136 344 137 345
rect 137 344 138 345
rect 138 344 139 345
rect 139 344 140 345
rect 510 344 511 345
rect 511 344 512 345
rect 512 344 513 345
rect 513 344 514 345
rect 514 344 515 345
rect 515 344 516 345
rect 516 344 517 345
rect 517 344 518 345
rect 518 344 519 345
rect 519 344 520 345
rect 520 344 521 345
rect 521 344 522 345
rect 522 344 523 345
rect 523 344 524 345
rect 524 344 525 345
rect 525 344 526 345
rect 526 344 527 345
rect 527 344 528 345
rect 528 344 529 345
rect 529 344 530 345
rect 530 344 531 345
rect 531 344 532 345
rect 532 344 533 345
rect 21 343 22 344
rect 22 343 23 344
rect 23 343 24 344
rect 24 343 25 344
rect 25 343 26 344
rect 26 343 27 344
rect 27 343 28 344
rect 28 343 29 344
rect 29 343 30 344
rect 30 343 31 344
rect 122 343 123 344
rect 123 343 124 344
rect 124 343 125 344
rect 125 343 126 344
rect 126 343 127 344
rect 127 343 128 344
rect 128 343 129 344
rect 129 343 130 344
rect 130 343 131 344
rect 131 343 132 344
rect 132 343 133 344
rect 133 343 134 344
rect 134 343 135 344
rect 135 343 136 344
rect 136 343 137 344
rect 137 343 138 344
rect 138 343 139 344
rect 139 343 140 344
rect 512 343 513 344
rect 513 343 514 344
rect 514 343 515 344
rect 515 343 516 344
rect 516 343 517 344
rect 517 343 518 344
rect 518 343 519 344
rect 519 343 520 344
rect 520 343 521 344
rect 521 343 522 344
rect 522 343 523 344
rect 523 343 524 344
rect 524 343 525 344
rect 525 343 526 344
rect 526 343 527 344
rect 527 343 528 344
rect 528 343 529 344
rect 529 343 530 344
rect 530 343 531 344
rect 531 343 532 344
rect 532 343 533 344
rect 21 342 22 343
rect 22 342 23 343
rect 23 342 24 343
rect 24 342 25 343
rect 25 342 26 343
rect 26 342 27 343
rect 27 342 28 343
rect 28 342 29 343
rect 29 342 30 343
rect 30 342 31 343
rect 120 342 121 343
rect 121 342 122 343
rect 122 342 123 343
rect 123 342 124 343
rect 124 342 125 343
rect 125 342 126 343
rect 126 342 127 343
rect 127 342 128 343
rect 128 342 129 343
rect 129 342 130 343
rect 130 342 131 343
rect 131 342 132 343
rect 132 342 133 343
rect 133 342 134 343
rect 134 342 135 343
rect 135 342 136 343
rect 136 342 137 343
rect 137 342 138 343
rect 138 342 139 343
rect 139 342 140 343
rect 512 342 513 343
rect 513 342 514 343
rect 514 342 515 343
rect 515 342 516 343
rect 516 342 517 343
rect 517 342 518 343
rect 518 342 519 343
rect 519 342 520 343
rect 520 342 521 343
rect 521 342 522 343
rect 522 342 523 343
rect 523 342 524 343
rect 524 342 525 343
rect 525 342 526 343
rect 526 342 527 343
rect 527 342 528 343
rect 528 342 529 343
rect 529 342 530 343
rect 530 342 531 343
rect 531 342 532 343
rect 532 342 533 343
rect 21 341 22 342
rect 22 341 23 342
rect 23 341 24 342
rect 24 341 25 342
rect 25 341 26 342
rect 26 341 27 342
rect 27 341 28 342
rect 28 341 29 342
rect 29 341 30 342
rect 30 341 31 342
rect 120 341 121 342
rect 121 341 122 342
rect 122 341 123 342
rect 123 341 124 342
rect 124 341 125 342
rect 125 341 126 342
rect 126 341 127 342
rect 127 341 128 342
rect 128 341 129 342
rect 129 341 130 342
rect 130 341 131 342
rect 131 341 132 342
rect 132 341 133 342
rect 133 341 134 342
rect 134 341 135 342
rect 135 341 136 342
rect 136 341 137 342
rect 137 341 138 342
rect 512 341 513 342
rect 513 341 514 342
rect 514 341 515 342
rect 515 341 516 342
rect 516 341 517 342
rect 517 341 518 342
rect 518 341 519 342
rect 519 341 520 342
rect 520 341 521 342
rect 521 341 522 342
rect 522 341 523 342
rect 523 341 524 342
rect 524 341 525 342
rect 525 341 526 342
rect 526 341 527 342
rect 527 341 528 342
rect 528 341 529 342
rect 529 341 530 342
rect 530 341 531 342
rect 531 341 532 342
rect 532 341 533 342
rect 21 340 22 341
rect 22 340 23 341
rect 23 340 24 341
rect 24 340 25 341
rect 25 340 26 341
rect 26 340 27 341
rect 27 340 28 341
rect 28 340 29 341
rect 29 340 30 341
rect 30 340 31 341
rect 31 340 32 341
rect 32 340 33 341
rect 118 340 119 341
rect 119 340 120 341
rect 120 340 121 341
rect 121 340 122 341
rect 122 340 123 341
rect 123 340 124 341
rect 124 340 125 341
rect 125 340 126 341
rect 126 340 127 341
rect 127 340 128 341
rect 128 340 129 341
rect 129 340 130 341
rect 130 340 131 341
rect 131 340 132 341
rect 132 340 133 341
rect 133 340 134 341
rect 134 340 135 341
rect 135 340 136 341
rect 136 340 137 341
rect 137 340 138 341
rect 512 340 513 341
rect 513 340 514 341
rect 514 340 515 341
rect 515 340 516 341
rect 516 340 517 341
rect 517 340 518 341
rect 518 340 519 341
rect 519 340 520 341
rect 520 340 521 341
rect 521 340 522 341
rect 522 340 523 341
rect 523 340 524 341
rect 524 340 525 341
rect 525 340 526 341
rect 526 340 527 341
rect 527 340 528 341
rect 528 340 529 341
rect 529 340 530 341
rect 530 340 531 341
rect 531 340 532 341
rect 532 340 533 341
rect 21 339 22 340
rect 22 339 23 340
rect 23 339 24 340
rect 24 339 25 340
rect 25 339 26 340
rect 26 339 27 340
rect 27 339 28 340
rect 28 339 29 340
rect 29 339 30 340
rect 30 339 31 340
rect 31 339 32 340
rect 32 339 33 340
rect 118 339 119 340
rect 119 339 120 340
rect 120 339 121 340
rect 121 339 122 340
rect 122 339 123 340
rect 123 339 124 340
rect 124 339 125 340
rect 125 339 126 340
rect 126 339 127 340
rect 127 339 128 340
rect 128 339 129 340
rect 129 339 130 340
rect 130 339 131 340
rect 131 339 132 340
rect 132 339 133 340
rect 133 339 134 340
rect 134 339 135 340
rect 135 339 136 340
rect 514 339 515 340
rect 515 339 516 340
rect 516 339 517 340
rect 517 339 518 340
rect 518 339 519 340
rect 519 339 520 340
rect 520 339 521 340
rect 521 339 522 340
rect 522 339 523 340
rect 523 339 524 340
rect 524 339 525 340
rect 525 339 526 340
rect 526 339 527 340
rect 527 339 528 340
rect 528 339 529 340
rect 529 339 530 340
rect 530 339 531 340
rect 531 339 532 340
rect 532 339 533 340
rect 21 338 22 339
rect 22 338 23 339
rect 23 338 24 339
rect 24 338 25 339
rect 25 338 26 339
rect 26 338 27 339
rect 27 338 28 339
rect 28 338 29 339
rect 29 338 30 339
rect 30 338 31 339
rect 31 338 32 339
rect 32 338 33 339
rect 118 338 119 339
rect 119 338 120 339
rect 120 338 121 339
rect 121 338 122 339
rect 122 338 123 339
rect 123 338 124 339
rect 124 338 125 339
rect 125 338 126 339
rect 126 338 127 339
rect 127 338 128 339
rect 128 338 129 339
rect 129 338 130 339
rect 130 338 131 339
rect 131 338 132 339
rect 132 338 133 339
rect 133 338 134 339
rect 134 338 135 339
rect 135 338 136 339
rect 514 338 515 339
rect 515 338 516 339
rect 516 338 517 339
rect 517 338 518 339
rect 518 338 519 339
rect 519 338 520 339
rect 520 338 521 339
rect 521 338 522 339
rect 522 338 523 339
rect 523 338 524 339
rect 524 338 525 339
rect 525 338 526 339
rect 526 338 527 339
rect 527 338 528 339
rect 528 338 529 339
rect 529 338 530 339
rect 530 338 531 339
rect 531 338 532 339
rect 532 338 533 339
rect 533 338 534 339
rect 534 338 535 339
rect 21 337 22 338
rect 22 337 23 338
rect 23 337 24 338
rect 24 337 25 338
rect 25 337 26 338
rect 26 337 27 338
rect 27 337 28 338
rect 28 337 29 338
rect 29 337 30 338
rect 30 337 31 338
rect 31 337 32 338
rect 32 337 33 338
rect 118 337 119 338
rect 119 337 120 338
rect 120 337 121 338
rect 121 337 122 338
rect 122 337 123 338
rect 123 337 124 338
rect 124 337 125 338
rect 125 337 126 338
rect 126 337 127 338
rect 127 337 128 338
rect 128 337 129 338
rect 129 337 130 338
rect 130 337 131 338
rect 131 337 132 338
rect 132 337 133 338
rect 133 337 134 338
rect 515 337 516 338
rect 516 337 517 338
rect 517 337 518 338
rect 518 337 519 338
rect 519 337 520 338
rect 520 337 521 338
rect 521 337 522 338
rect 522 337 523 338
rect 523 337 524 338
rect 524 337 525 338
rect 525 337 526 338
rect 526 337 527 338
rect 527 337 528 338
rect 528 337 529 338
rect 529 337 530 338
rect 530 337 531 338
rect 531 337 532 338
rect 532 337 533 338
rect 533 337 534 338
rect 534 337 535 338
rect 21 336 22 337
rect 22 336 23 337
rect 23 336 24 337
rect 24 336 25 337
rect 25 336 26 337
rect 26 336 27 337
rect 27 336 28 337
rect 28 336 29 337
rect 29 336 30 337
rect 30 336 31 337
rect 31 336 32 337
rect 32 336 33 337
rect 33 336 34 337
rect 34 336 35 337
rect 117 336 118 337
rect 118 336 119 337
rect 119 336 120 337
rect 120 336 121 337
rect 121 336 122 337
rect 122 336 123 337
rect 123 336 124 337
rect 124 336 125 337
rect 125 336 126 337
rect 126 336 127 337
rect 127 336 128 337
rect 128 336 129 337
rect 129 336 130 337
rect 130 336 131 337
rect 131 336 132 337
rect 132 336 133 337
rect 133 336 134 337
rect 515 336 516 337
rect 516 336 517 337
rect 517 336 518 337
rect 518 336 519 337
rect 519 336 520 337
rect 520 336 521 337
rect 521 336 522 337
rect 522 336 523 337
rect 523 336 524 337
rect 524 336 525 337
rect 525 336 526 337
rect 526 336 527 337
rect 527 336 528 337
rect 528 336 529 337
rect 529 336 530 337
rect 530 336 531 337
rect 531 336 532 337
rect 532 336 533 337
rect 533 336 534 337
rect 534 336 535 337
rect 21 335 22 336
rect 22 335 23 336
rect 23 335 24 336
rect 24 335 25 336
rect 25 335 26 336
rect 26 335 27 336
rect 27 335 28 336
rect 28 335 29 336
rect 29 335 30 336
rect 30 335 31 336
rect 31 335 32 336
rect 32 335 33 336
rect 33 335 34 336
rect 34 335 35 336
rect 117 335 118 336
rect 118 335 119 336
rect 119 335 120 336
rect 120 335 121 336
rect 121 335 122 336
rect 122 335 123 336
rect 123 335 124 336
rect 124 335 125 336
rect 125 335 126 336
rect 126 335 127 336
rect 127 335 128 336
rect 128 335 129 336
rect 129 335 130 336
rect 130 335 131 336
rect 131 335 132 336
rect 132 335 133 336
rect 515 335 516 336
rect 516 335 517 336
rect 517 335 518 336
rect 518 335 519 336
rect 519 335 520 336
rect 520 335 521 336
rect 521 335 522 336
rect 522 335 523 336
rect 523 335 524 336
rect 524 335 525 336
rect 525 335 526 336
rect 526 335 527 336
rect 527 335 528 336
rect 528 335 529 336
rect 529 335 530 336
rect 530 335 531 336
rect 531 335 532 336
rect 532 335 533 336
rect 533 335 534 336
rect 534 335 535 336
rect 21 334 22 335
rect 22 334 23 335
rect 23 334 24 335
rect 24 334 25 335
rect 25 334 26 335
rect 26 334 27 335
rect 27 334 28 335
rect 28 334 29 335
rect 29 334 30 335
rect 30 334 31 335
rect 31 334 32 335
rect 32 334 33 335
rect 33 334 34 335
rect 34 334 35 335
rect 117 334 118 335
rect 118 334 119 335
rect 119 334 120 335
rect 120 334 121 335
rect 121 334 122 335
rect 122 334 123 335
rect 123 334 124 335
rect 124 334 125 335
rect 125 334 126 335
rect 126 334 127 335
rect 127 334 128 335
rect 128 334 129 335
rect 129 334 130 335
rect 130 334 131 335
rect 131 334 132 335
rect 132 334 133 335
rect 515 334 516 335
rect 516 334 517 335
rect 517 334 518 335
rect 518 334 519 335
rect 519 334 520 335
rect 520 334 521 335
rect 521 334 522 335
rect 522 334 523 335
rect 523 334 524 335
rect 524 334 525 335
rect 525 334 526 335
rect 526 334 527 335
rect 527 334 528 335
rect 528 334 529 335
rect 529 334 530 335
rect 530 334 531 335
rect 531 334 532 335
rect 532 334 533 335
rect 533 334 534 335
rect 534 334 535 335
rect 21 333 22 334
rect 22 333 23 334
rect 23 333 24 334
rect 24 333 25 334
rect 25 333 26 334
rect 26 333 27 334
rect 27 333 28 334
rect 28 333 29 334
rect 29 333 30 334
rect 30 333 31 334
rect 31 333 32 334
rect 32 333 33 334
rect 33 333 34 334
rect 34 333 35 334
rect 117 333 118 334
rect 118 333 119 334
rect 119 333 120 334
rect 120 333 121 334
rect 121 333 122 334
rect 122 333 123 334
rect 123 333 124 334
rect 124 333 125 334
rect 125 333 126 334
rect 126 333 127 334
rect 127 333 128 334
rect 128 333 129 334
rect 129 333 130 334
rect 130 333 131 334
rect 517 333 518 334
rect 518 333 519 334
rect 519 333 520 334
rect 520 333 521 334
rect 521 333 522 334
rect 522 333 523 334
rect 523 333 524 334
rect 524 333 525 334
rect 525 333 526 334
rect 526 333 527 334
rect 527 333 528 334
rect 528 333 529 334
rect 529 333 530 334
rect 530 333 531 334
rect 531 333 532 334
rect 532 333 533 334
rect 533 333 534 334
rect 534 333 535 334
rect 21 332 22 333
rect 22 332 23 333
rect 23 332 24 333
rect 24 332 25 333
rect 25 332 26 333
rect 26 332 27 333
rect 27 332 28 333
rect 28 332 29 333
rect 29 332 30 333
rect 30 332 31 333
rect 31 332 32 333
rect 32 332 33 333
rect 33 332 34 333
rect 34 332 35 333
rect 35 332 36 333
rect 36 332 37 333
rect 115 332 116 333
rect 116 332 117 333
rect 117 332 118 333
rect 118 332 119 333
rect 119 332 120 333
rect 120 332 121 333
rect 121 332 122 333
rect 122 332 123 333
rect 123 332 124 333
rect 124 332 125 333
rect 125 332 126 333
rect 126 332 127 333
rect 127 332 128 333
rect 128 332 129 333
rect 129 332 130 333
rect 130 332 131 333
rect 517 332 518 333
rect 518 332 519 333
rect 519 332 520 333
rect 520 332 521 333
rect 521 332 522 333
rect 522 332 523 333
rect 523 332 524 333
rect 524 332 525 333
rect 525 332 526 333
rect 526 332 527 333
rect 527 332 528 333
rect 528 332 529 333
rect 529 332 530 333
rect 530 332 531 333
rect 531 332 532 333
rect 532 332 533 333
rect 533 332 534 333
rect 534 332 535 333
rect 21 331 22 332
rect 22 331 23 332
rect 23 331 24 332
rect 24 331 25 332
rect 25 331 26 332
rect 26 331 27 332
rect 27 331 28 332
rect 28 331 29 332
rect 29 331 30 332
rect 30 331 31 332
rect 31 331 32 332
rect 32 331 33 332
rect 33 331 34 332
rect 34 331 35 332
rect 35 331 36 332
rect 36 331 37 332
rect 115 331 116 332
rect 116 331 117 332
rect 117 331 118 332
rect 118 331 119 332
rect 119 331 120 332
rect 120 331 121 332
rect 121 331 122 332
rect 122 331 123 332
rect 123 331 124 332
rect 124 331 125 332
rect 125 331 126 332
rect 126 331 127 332
rect 127 331 128 332
rect 128 331 129 332
rect 517 331 518 332
rect 518 331 519 332
rect 519 331 520 332
rect 520 331 521 332
rect 521 331 522 332
rect 522 331 523 332
rect 523 331 524 332
rect 524 331 525 332
rect 525 331 526 332
rect 526 331 527 332
rect 527 331 528 332
rect 528 331 529 332
rect 529 331 530 332
rect 530 331 531 332
rect 531 331 532 332
rect 532 331 533 332
rect 533 331 534 332
rect 534 331 535 332
rect 21 330 22 331
rect 22 330 23 331
rect 23 330 24 331
rect 24 330 25 331
rect 25 330 26 331
rect 26 330 27 331
rect 27 330 28 331
rect 28 330 29 331
rect 29 330 30 331
rect 30 330 31 331
rect 31 330 32 331
rect 32 330 33 331
rect 33 330 34 331
rect 34 330 35 331
rect 35 330 36 331
rect 36 330 37 331
rect 115 330 116 331
rect 116 330 117 331
rect 117 330 118 331
rect 118 330 119 331
rect 119 330 120 331
rect 120 330 121 331
rect 121 330 122 331
rect 122 330 123 331
rect 123 330 124 331
rect 124 330 125 331
rect 125 330 126 331
rect 126 330 127 331
rect 127 330 128 331
rect 128 330 129 331
rect 517 330 518 331
rect 518 330 519 331
rect 519 330 520 331
rect 520 330 521 331
rect 521 330 522 331
rect 522 330 523 331
rect 523 330 524 331
rect 524 330 525 331
rect 525 330 526 331
rect 526 330 527 331
rect 527 330 528 331
rect 528 330 529 331
rect 529 330 530 331
rect 530 330 531 331
rect 531 330 532 331
rect 532 330 533 331
rect 533 330 534 331
rect 534 330 535 331
rect 21 329 22 330
rect 22 329 23 330
rect 23 329 24 330
rect 24 329 25 330
rect 25 329 26 330
rect 26 329 27 330
rect 27 329 28 330
rect 28 329 29 330
rect 29 329 30 330
rect 30 329 31 330
rect 31 329 32 330
rect 32 329 33 330
rect 33 329 34 330
rect 34 329 35 330
rect 35 329 36 330
rect 36 329 37 330
rect 115 329 116 330
rect 116 329 117 330
rect 117 329 118 330
rect 118 329 119 330
rect 119 329 120 330
rect 120 329 121 330
rect 121 329 122 330
rect 122 329 123 330
rect 123 329 124 330
rect 124 329 125 330
rect 125 329 126 330
rect 126 329 127 330
rect 127 329 128 330
rect 128 329 129 330
rect 517 329 518 330
rect 518 329 519 330
rect 519 329 520 330
rect 520 329 521 330
rect 521 329 522 330
rect 522 329 523 330
rect 523 329 524 330
rect 524 329 525 330
rect 525 329 526 330
rect 526 329 527 330
rect 527 329 528 330
rect 528 329 529 330
rect 529 329 530 330
rect 530 329 531 330
rect 531 329 532 330
rect 532 329 533 330
rect 533 329 534 330
rect 534 329 535 330
rect 21 328 22 329
rect 22 328 23 329
rect 23 328 24 329
rect 24 328 25 329
rect 25 328 26 329
rect 26 328 27 329
rect 27 328 28 329
rect 28 328 29 329
rect 29 328 30 329
rect 30 328 31 329
rect 31 328 32 329
rect 32 328 33 329
rect 33 328 34 329
rect 34 328 35 329
rect 35 328 36 329
rect 36 328 37 329
rect 115 328 116 329
rect 116 328 117 329
rect 117 328 118 329
rect 118 328 119 329
rect 119 328 120 329
rect 120 328 121 329
rect 121 328 122 329
rect 122 328 123 329
rect 123 328 124 329
rect 124 328 125 329
rect 125 328 126 329
rect 126 328 127 329
rect 519 328 520 329
rect 520 328 521 329
rect 521 328 522 329
rect 522 328 523 329
rect 523 328 524 329
rect 524 328 525 329
rect 525 328 526 329
rect 526 328 527 329
rect 527 328 528 329
rect 528 328 529 329
rect 529 328 530 329
rect 530 328 531 329
rect 531 328 532 329
rect 532 328 533 329
rect 533 328 534 329
rect 534 328 535 329
rect 21 327 22 328
rect 22 327 23 328
rect 23 327 24 328
rect 24 327 25 328
rect 25 327 26 328
rect 26 327 27 328
rect 27 327 28 328
rect 28 327 29 328
rect 29 327 30 328
rect 30 327 31 328
rect 31 327 32 328
rect 32 327 33 328
rect 33 327 34 328
rect 34 327 35 328
rect 35 327 36 328
rect 36 327 37 328
rect 37 327 38 328
rect 38 327 39 328
rect 113 327 114 328
rect 114 327 115 328
rect 115 327 116 328
rect 116 327 117 328
rect 117 327 118 328
rect 118 327 119 328
rect 119 327 120 328
rect 120 327 121 328
rect 121 327 122 328
rect 122 327 123 328
rect 123 327 124 328
rect 124 327 125 328
rect 125 327 126 328
rect 126 327 127 328
rect 519 327 520 328
rect 520 327 521 328
rect 521 327 522 328
rect 522 327 523 328
rect 523 327 524 328
rect 524 327 525 328
rect 525 327 526 328
rect 526 327 527 328
rect 527 327 528 328
rect 528 327 529 328
rect 529 327 530 328
rect 530 327 531 328
rect 531 327 532 328
rect 532 327 533 328
rect 533 327 534 328
rect 534 327 535 328
rect 535 327 536 328
rect 536 327 537 328
rect 21 326 22 327
rect 22 326 23 327
rect 23 326 24 327
rect 24 326 25 327
rect 25 326 26 327
rect 26 326 27 327
rect 27 326 28 327
rect 28 326 29 327
rect 29 326 30 327
rect 30 326 31 327
rect 31 326 32 327
rect 32 326 33 327
rect 33 326 34 327
rect 34 326 35 327
rect 35 326 36 327
rect 36 326 37 327
rect 37 326 38 327
rect 38 326 39 327
rect 113 326 114 327
rect 114 326 115 327
rect 115 326 116 327
rect 116 326 117 327
rect 117 326 118 327
rect 118 326 119 327
rect 119 326 120 327
rect 120 326 121 327
rect 121 326 122 327
rect 122 326 123 327
rect 123 326 124 327
rect 124 326 125 327
rect 125 326 126 327
rect 126 326 127 327
rect 521 326 522 327
rect 522 326 523 327
rect 523 326 524 327
rect 524 326 525 327
rect 525 326 526 327
rect 526 326 527 327
rect 527 326 528 327
rect 528 326 529 327
rect 529 326 530 327
rect 530 326 531 327
rect 531 326 532 327
rect 532 326 533 327
rect 533 326 534 327
rect 534 326 535 327
rect 535 326 536 327
rect 536 326 537 327
rect 21 325 22 326
rect 22 325 23 326
rect 23 325 24 326
rect 24 325 25 326
rect 25 325 26 326
rect 26 325 27 326
rect 27 325 28 326
rect 28 325 29 326
rect 29 325 30 326
rect 30 325 31 326
rect 31 325 32 326
rect 32 325 33 326
rect 33 325 34 326
rect 34 325 35 326
rect 35 325 36 326
rect 36 325 37 326
rect 37 325 38 326
rect 38 325 39 326
rect 39 325 40 326
rect 40 325 41 326
rect 113 325 114 326
rect 114 325 115 326
rect 115 325 116 326
rect 116 325 117 326
rect 117 325 118 326
rect 118 325 119 326
rect 119 325 120 326
rect 120 325 121 326
rect 121 325 122 326
rect 122 325 123 326
rect 123 325 124 326
rect 124 325 125 326
rect 125 325 126 326
rect 126 325 127 326
rect 521 325 522 326
rect 522 325 523 326
rect 523 325 524 326
rect 524 325 525 326
rect 525 325 526 326
rect 526 325 527 326
rect 527 325 528 326
rect 528 325 529 326
rect 529 325 530 326
rect 530 325 531 326
rect 531 325 532 326
rect 532 325 533 326
rect 533 325 534 326
rect 534 325 535 326
rect 535 325 536 326
rect 536 325 537 326
rect 23 324 24 325
rect 24 324 25 325
rect 25 324 26 325
rect 26 324 27 325
rect 27 324 28 325
rect 28 324 29 325
rect 29 324 30 325
rect 30 324 31 325
rect 31 324 32 325
rect 32 324 33 325
rect 33 324 34 325
rect 34 324 35 325
rect 35 324 36 325
rect 36 324 37 325
rect 37 324 38 325
rect 38 324 39 325
rect 39 324 40 325
rect 40 324 41 325
rect 113 324 114 325
rect 114 324 115 325
rect 115 324 116 325
rect 116 324 117 325
rect 117 324 118 325
rect 118 324 119 325
rect 119 324 120 325
rect 120 324 121 325
rect 121 324 122 325
rect 122 324 123 325
rect 123 324 124 325
rect 124 324 125 325
rect 521 324 522 325
rect 522 324 523 325
rect 523 324 524 325
rect 524 324 525 325
rect 525 324 526 325
rect 526 324 527 325
rect 527 324 528 325
rect 528 324 529 325
rect 529 324 530 325
rect 530 324 531 325
rect 531 324 532 325
rect 532 324 533 325
rect 533 324 534 325
rect 534 324 535 325
rect 535 324 536 325
rect 536 324 537 325
rect 23 323 24 324
rect 24 323 25 324
rect 25 323 26 324
rect 26 323 27 324
rect 27 323 28 324
rect 28 323 29 324
rect 29 323 30 324
rect 30 323 31 324
rect 31 323 32 324
rect 32 323 33 324
rect 33 323 34 324
rect 34 323 35 324
rect 35 323 36 324
rect 36 323 37 324
rect 37 323 38 324
rect 38 323 39 324
rect 39 323 40 324
rect 40 323 41 324
rect 111 323 112 324
rect 112 323 113 324
rect 113 323 114 324
rect 114 323 115 324
rect 115 323 116 324
rect 116 323 117 324
rect 117 323 118 324
rect 118 323 119 324
rect 119 323 120 324
rect 120 323 121 324
rect 121 323 122 324
rect 122 323 123 324
rect 123 323 124 324
rect 124 323 125 324
rect 521 323 522 324
rect 522 323 523 324
rect 523 323 524 324
rect 524 323 525 324
rect 525 323 526 324
rect 526 323 527 324
rect 527 323 528 324
rect 528 323 529 324
rect 529 323 530 324
rect 530 323 531 324
rect 531 323 532 324
rect 532 323 533 324
rect 533 323 534 324
rect 534 323 535 324
rect 535 323 536 324
rect 536 323 537 324
rect 23 322 24 323
rect 24 322 25 323
rect 25 322 26 323
rect 26 322 27 323
rect 27 322 28 323
rect 28 322 29 323
rect 29 322 30 323
rect 30 322 31 323
rect 31 322 32 323
rect 32 322 33 323
rect 33 322 34 323
rect 34 322 35 323
rect 35 322 36 323
rect 36 322 37 323
rect 37 322 38 323
rect 38 322 39 323
rect 39 322 40 323
rect 40 322 41 323
rect 111 322 112 323
rect 112 322 113 323
rect 113 322 114 323
rect 114 322 115 323
rect 115 322 116 323
rect 116 322 117 323
rect 117 322 118 323
rect 118 322 119 323
rect 119 322 120 323
rect 120 322 121 323
rect 121 322 122 323
rect 122 322 123 323
rect 521 322 522 323
rect 522 322 523 323
rect 523 322 524 323
rect 524 322 525 323
rect 525 322 526 323
rect 526 322 527 323
rect 527 322 528 323
rect 528 322 529 323
rect 529 322 530 323
rect 530 322 531 323
rect 531 322 532 323
rect 532 322 533 323
rect 533 322 534 323
rect 534 322 535 323
rect 535 322 536 323
rect 536 322 537 323
rect 23 321 24 322
rect 24 321 25 322
rect 25 321 26 322
rect 26 321 27 322
rect 27 321 28 322
rect 28 321 29 322
rect 29 321 30 322
rect 30 321 31 322
rect 31 321 32 322
rect 32 321 33 322
rect 33 321 34 322
rect 34 321 35 322
rect 35 321 36 322
rect 36 321 37 322
rect 37 321 38 322
rect 38 321 39 322
rect 39 321 40 322
rect 40 321 41 322
rect 41 321 42 322
rect 42 321 43 322
rect 111 321 112 322
rect 112 321 113 322
rect 113 321 114 322
rect 114 321 115 322
rect 115 321 116 322
rect 116 321 117 322
rect 117 321 118 322
rect 118 321 119 322
rect 119 321 120 322
rect 120 321 121 322
rect 121 321 122 322
rect 122 321 123 322
rect 521 321 522 322
rect 522 321 523 322
rect 523 321 524 322
rect 524 321 525 322
rect 525 321 526 322
rect 526 321 527 322
rect 527 321 528 322
rect 528 321 529 322
rect 529 321 530 322
rect 530 321 531 322
rect 531 321 532 322
rect 532 321 533 322
rect 533 321 534 322
rect 534 321 535 322
rect 535 321 536 322
rect 536 321 537 322
rect 23 320 24 321
rect 24 320 25 321
rect 25 320 26 321
rect 26 320 27 321
rect 27 320 28 321
rect 28 320 29 321
rect 29 320 30 321
rect 30 320 31 321
rect 31 320 32 321
rect 32 320 33 321
rect 33 320 34 321
rect 34 320 35 321
rect 35 320 36 321
rect 36 320 37 321
rect 37 320 38 321
rect 38 320 39 321
rect 39 320 40 321
rect 40 320 41 321
rect 41 320 42 321
rect 42 320 43 321
rect 111 320 112 321
rect 112 320 113 321
rect 113 320 114 321
rect 114 320 115 321
rect 115 320 116 321
rect 116 320 117 321
rect 117 320 118 321
rect 118 320 119 321
rect 119 320 120 321
rect 120 320 121 321
rect 523 320 524 321
rect 524 320 525 321
rect 525 320 526 321
rect 526 320 527 321
rect 527 320 528 321
rect 528 320 529 321
rect 529 320 530 321
rect 530 320 531 321
rect 531 320 532 321
rect 532 320 533 321
rect 533 320 534 321
rect 534 320 535 321
rect 535 320 536 321
rect 536 320 537 321
rect 23 319 24 320
rect 24 319 25 320
rect 25 319 26 320
rect 26 319 27 320
rect 27 319 28 320
rect 28 319 29 320
rect 29 319 30 320
rect 30 319 31 320
rect 31 319 32 320
rect 32 319 33 320
rect 33 319 34 320
rect 34 319 35 320
rect 35 319 36 320
rect 36 319 37 320
rect 37 319 38 320
rect 38 319 39 320
rect 39 319 40 320
rect 40 319 41 320
rect 41 319 42 320
rect 42 319 43 320
rect 43 319 44 320
rect 44 319 45 320
rect 111 319 112 320
rect 112 319 113 320
rect 113 319 114 320
rect 114 319 115 320
rect 115 319 116 320
rect 116 319 117 320
rect 117 319 118 320
rect 118 319 119 320
rect 119 319 120 320
rect 120 319 121 320
rect 523 319 524 320
rect 524 319 525 320
rect 525 319 526 320
rect 526 319 527 320
rect 527 319 528 320
rect 528 319 529 320
rect 529 319 530 320
rect 530 319 531 320
rect 531 319 532 320
rect 532 319 533 320
rect 533 319 534 320
rect 534 319 535 320
rect 535 319 536 320
rect 536 319 537 320
rect 25 318 26 319
rect 26 318 27 319
rect 27 318 28 319
rect 28 318 29 319
rect 29 318 30 319
rect 30 318 31 319
rect 31 318 32 319
rect 32 318 33 319
rect 33 318 34 319
rect 34 318 35 319
rect 35 318 36 319
rect 36 318 37 319
rect 37 318 38 319
rect 38 318 39 319
rect 39 318 40 319
rect 40 318 41 319
rect 41 318 42 319
rect 42 318 43 319
rect 43 318 44 319
rect 44 318 45 319
rect 111 318 112 319
rect 112 318 113 319
rect 113 318 114 319
rect 114 318 115 319
rect 115 318 116 319
rect 116 318 117 319
rect 117 318 118 319
rect 118 318 119 319
rect 525 318 526 319
rect 526 318 527 319
rect 527 318 528 319
rect 528 318 529 319
rect 529 318 530 319
rect 530 318 531 319
rect 531 318 532 319
rect 532 318 533 319
rect 533 318 534 319
rect 534 318 535 319
rect 535 318 536 319
rect 536 318 537 319
rect 25 317 26 318
rect 26 317 27 318
rect 27 317 28 318
rect 28 317 29 318
rect 29 317 30 318
rect 30 317 31 318
rect 31 317 32 318
rect 32 317 33 318
rect 33 317 34 318
rect 34 317 35 318
rect 35 317 36 318
rect 36 317 37 318
rect 37 317 38 318
rect 38 317 39 318
rect 39 317 40 318
rect 40 317 41 318
rect 41 317 42 318
rect 42 317 43 318
rect 43 317 44 318
rect 44 317 45 318
rect 45 317 46 318
rect 109 317 110 318
rect 110 317 111 318
rect 111 317 112 318
rect 112 317 113 318
rect 113 317 114 318
rect 114 317 115 318
rect 115 317 116 318
rect 116 317 117 318
rect 117 317 118 318
rect 118 317 119 318
rect 525 317 526 318
rect 526 317 527 318
rect 527 317 528 318
rect 528 317 529 318
rect 529 317 530 318
rect 530 317 531 318
rect 531 317 532 318
rect 532 317 533 318
rect 533 317 534 318
rect 534 317 535 318
rect 535 317 536 318
rect 536 317 537 318
rect 25 316 26 317
rect 26 316 27 317
rect 27 316 28 317
rect 28 316 29 317
rect 29 316 30 317
rect 30 316 31 317
rect 31 316 32 317
rect 32 316 33 317
rect 33 316 34 317
rect 34 316 35 317
rect 35 316 36 317
rect 36 316 37 317
rect 37 316 38 317
rect 38 316 39 317
rect 39 316 40 317
rect 40 316 41 317
rect 41 316 42 317
rect 42 316 43 317
rect 43 316 44 317
rect 44 316 45 317
rect 45 316 46 317
rect 109 316 110 317
rect 110 316 111 317
rect 111 316 112 317
rect 112 316 113 317
rect 113 316 114 317
rect 114 316 115 317
rect 115 316 116 317
rect 116 316 117 317
rect 117 316 118 317
rect 118 316 119 317
rect 525 316 526 317
rect 526 316 527 317
rect 527 316 528 317
rect 528 316 529 317
rect 529 316 530 317
rect 530 316 531 317
rect 531 316 532 317
rect 532 316 533 317
rect 533 316 534 317
rect 534 316 535 317
rect 535 316 536 317
rect 536 316 537 317
rect 25 315 26 316
rect 26 315 27 316
rect 27 315 28 316
rect 28 315 29 316
rect 29 315 30 316
rect 30 315 31 316
rect 31 315 32 316
rect 32 315 33 316
rect 33 315 34 316
rect 34 315 35 316
rect 35 315 36 316
rect 36 315 37 316
rect 37 315 38 316
rect 38 315 39 316
rect 39 315 40 316
rect 40 315 41 316
rect 41 315 42 316
rect 42 315 43 316
rect 43 315 44 316
rect 44 315 45 316
rect 45 315 46 316
rect 109 315 110 316
rect 110 315 111 316
rect 111 315 112 316
rect 112 315 113 316
rect 113 315 114 316
rect 114 315 115 316
rect 115 315 116 316
rect 116 315 117 316
rect 117 315 118 316
rect 118 315 119 316
rect 525 315 526 316
rect 526 315 527 316
rect 527 315 528 316
rect 528 315 529 316
rect 529 315 530 316
rect 530 315 531 316
rect 531 315 532 316
rect 532 315 533 316
rect 533 315 534 316
rect 534 315 535 316
rect 535 315 536 316
rect 536 315 537 316
rect 27 314 28 315
rect 28 314 29 315
rect 29 314 30 315
rect 30 314 31 315
rect 31 314 32 315
rect 32 314 33 315
rect 33 314 34 315
rect 34 314 35 315
rect 35 314 36 315
rect 36 314 37 315
rect 37 314 38 315
rect 38 314 39 315
rect 39 314 40 315
rect 40 314 41 315
rect 41 314 42 315
rect 42 314 43 315
rect 43 314 44 315
rect 44 314 45 315
rect 45 314 46 315
rect 109 314 110 315
rect 110 314 111 315
rect 111 314 112 315
rect 112 314 113 315
rect 113 314 114 315
rect 114 314 115 315
rect 115 314 116 315
rect 116 314 117 315
rect 117 314 118 315
rect 525 314 526 315
rect 526 314 527 315
rect 527 314 528 315
rect 528 314 529 315
rect 529 314 530 315
rect 530 314 531 315
rect 531 314 532 315
rect 532 314 533 315
rect 533 314 534 315
rect 534 314 535 315
rect 535 314 536 315
rect 536 314 537 315
rect 27 313 28 314
rect 28 313 29 314
rect 29 313 30 314
rect 30 313 31 314
rect 31 313 32 314
rect 32 313 33 314
rect 33 313 34 314
rect 34 313 35 314
rect 35 313 36 314
rect 36 313 37 314
rect 37 313 38 314
rect 38 313 39 314
rect 39 313 40 314
rect 40 313 41 314
rect 41 313 42 314
rect 42 313 43 314
rect 43 313 44 314
rect 44 313 45 314
rect 45 313 46 314
rect 46 313 47 314
rect 47 313 48 314
rect 107 313 108 314
rect 108 313 109 314
rect 109 313 110 314
rect 110 313 111 314
rect 111 313 112 314
rect 112 313 113 314
rect 113 313 114 314
rect 114 313 115 314
rect 115 313 116 314
rect 116 313 117 314
rect 117 313 118 314
rect 525 313 526 314
rect 526 313 527 314
rect 527 313 528 314
rect 528 313 529 314
rect 529 313 530 314
rect 530 313 531 314
rect 531 313 532 314
rect 532 313 533 314
rect 533 313 534 314
rect 534 313 535 314
rect 535 313 536 314
rect 536 313 537 314
rect 29 312 30 313
rect 30 312 31 313
rect 31 312 32 313
rect 32 312 33 313
rect 33 312 34 313
rect 34 312 35 313
rect 35 312 36 313
rect 36 312 37 313
rect 37 312 38 313
rect 38 312 39 313
rect 39 312 40 313
rect 40 312 41 313
rect 41 312 42 313
rect 42 312 43 313
rect 43 312 44 313
rect 44 312 45 313
rect 45 312 46 313
rect 46 312 47 313
rect 47 312 48 313
rect 107 312 108 313
rect 108 312 109 313
rect 109 312 110 313
rect 110 312 111 313
rect 111 312 112 313
rect 112 312 113 313
rect 113 312 114 313
rect 114 312 115 313
rect 115 312 116 313
rect 525 312 526 313
rect 526 312 527 313
rect 527 312 528 313
rect 528 312 529 313
rect 529 312 530 313
rect 530 312 531 313
rect 531 312 532 313
rect 532 312 533 313
rect 533 312 534 313
rect 534 312 535 313
rect 535 312 536 313
rect 536 312 537 313
rect 29 311 30 312
rect 30 311 31 312
rect 31 311 32 312
rect 32 311 33 312
rect 33 311 34 312
rect 34 311 35 312
rect 35 311 36 312
rect 36 311 37 312
rect 37 311 38 312
rect 38 311 39 312
rect 39 311 40 312
rect 40 311 41 312
rect 41 311 42 312
rect 42 311 43 312
rect 43 311 44 312
rect 44 311 45 312
rect 45 311 46 312
rect 46 311 47 312
rect 47 311 48 312
rect 48 311 49 312
rect 49 311 50 312
rect 107 311 108 312
rect 108 311 109 312
rect 109 311 110 312
rect 110 311 111 312
rect 111 311 112 312
rect 112 311 113 312
rect 113 311 114 312
rect 114 311 115 312
rect 115 311 116 312
rect 525 311 526 312
rect 526 311 527 312
rect 527 311 528 312
rect 528 311 529 312
rect 529 311 530 312
rect 530 311 531 312
rect 531 311 532 312
rect 532 311 533 312
rect 533 311 534 312
rect 534 311 535 312
rect 535 311 536 312
rect 536 311 537 312
rect 537 311 538 312
rect 538 311 539 312
rect 29 310 30 311
rect 30 310 31 311
rect 31 310 32 311
rect 32 310 33 311
rect 33 310 34 311
rect 34 310 35 311
rect 35 310 36 311
rect 36 310 37 311
rect 37 310 38 311
rect 38 310 39 311
rect 39 310 40 311
rect 40 310 41 311
rect 41 310 42 311
rect 42 310 43 311
rect 43 310 44 311
rect 44 310 45 311
rect 45 310 46 311
rect 46 310 47 311
rect 47 310 48 311
rect 48 310 49 311
rect 49 310 50 311
rect 107 310 108 311
rect 108 310 109 311
rect 109 310 110 311
rect 110 310 111 311
rect 111 310 112 311
rect 112 310 113 311
rect 113 310 114 311
rect 114 310 115 311
rect 115 310 116 311
rect 527 310 528 311
rect 528 310 529 311
rect 529 310 530 311
rect 530 310 531 311
rect 531 310 532 311
rect 532 310 533 311
rect 533 310 534 311
rect 534 310 535 311
rect 535 310 536 311
rect 536 310 537 311
rect 537 310 538 311
rect 538 310 539 311
rect 29 309 30 310
rect 30 309 31 310
rect 31 309 32 310
rect 32 309 33 310
rect 33 309 34 310
rect 34 309 35 310
rect 35 309 36 310
rect 36 309 37 310
rect 37 309 38 310
rect 38 309 39 310
rect 39 309 40 310
rect 40 309 41 310
rect 41 309 42 310
rect 42 309 43 310
rect 43 309 44 310
rect 44 309 45 310
rect 45 309 46 310
rect 46 309 47 310
rect 47 309 48 310
rect 48 309 49 310
rect 49 309 50 310
rect 50 309 51 310
rect 51 309 52 310
rect 105 309 106 310
rect 106 309 107 310
rect 107 309 108 310
rect 108 309 109 310
rect 109 309 110 310
rect 110 309 111 310
rect 111 309 112 310
rect 112 309 113 310
rect 113 309 114 310
rect 114 309 115 310
rect 115 309 116 310
rect 527 309 528 310
rect 528 309 529 310
rect 529 309 530 310
rect 530 309 531 310
rect 531 309 532 310
rect 532 309 533 310
rect 533 309 534 310
rect 534 309 535 310
rect 535 309 536 310
rect 536 309 537 310
rect 537 309 538 310
rect 538 309 539 310
rect 32 308 33 309
rect 33 308 34 309
rect 34 308 35 309
rect 35 308 36 309
rect 36 308 37 309
rect 37 308 38 309
rect 38 308 39 309
rect 39 308 40 309
rect 40 308 41 309
rect 41 308 42 309
rect 42 308 43 309
rect 43 308 44 309
rect 44 308 45 309
rect 45 308 46 309
rect 46 308 47 309
rect 47 308 48 309
rect 48 308 49 309
rect 49 308 50 309
rect 50 308 51 309
rect 51 308 52 309
rect 105 308 106 309
rect 106 308 107 309
rect 107 308 108 309
rect 108 308 109 309
rect 109 308 110 309
rect 110 308 111 309
rect 111 308 112 309
rect 112 308 113 309
rect 113 308 114 309
rect 527 308 528 309
rect 528 308 529 309
rect 529 308 530 309
rect 530 308 531 309
rect 531 308 532 309
rect 532 308 533 309
rect 533 308 534 309
rect 534 308 535 309
rect 535 308 536 309
rect 536 308 537 309
rect 537 308 538 309
rect 538 308 539 309
rect 32 307 33 308
rect 33 307 34 308
rect 34 307 35 308
rect 35 307 36 308
rect 36 307 37 308
rect 37 307 38 308
rect 38 307 39 308
rect 39 307 40 308
rect 40 307 41 308
rect 41 307 42 308
rect 42 307 43 308
rect 43 307 44 308
rect 44 307 45 308
rect 45 307 46 308
rect 46 307 47 308
rect 47 307 48 308
rect 48 307 49 308
rect 49 307 50 308
rect 50 307 51 308
rect 51 307 52 308
rect 52 307 53 308
rect 53 307 54 308
rect 54 307 55 308
rect 55 307 56 308
rect 105 307 106 308
rect 106 307 107 308
rect 107 307 108 308
rect 108 307 109 308
rect 109 307 110 308
rect 110 307 111 308
rect 111 307 112 308
rect 112 307 113 308
rect 113 307 114 308
rect 527 307 528 308
rect 528 307 529 308
rect 529 307 530 308
rect 530 307 531 308
rect 531 307 532 308
rect 532 307 533 308
rect 533 307 534 308
rect 534 307 535 308
rect 535 307 536 308
rect 536 307 537 308
rect 537 307 538 308
rect 538 307 539 308
rect 34 306 35 307
rect 35 306 36 307
rect 36 306 37 307
rect 37 306 38 307
rect 38 306 39 307
rect 39 306 40 307
rect 40 306 41 307
rect 41 306 42 307
rect 42 306 43 307
rect 43 306 44 307
rect 44 306 45 307
rect 45 306 46 307
rect 46 306 47 307
rect 47 306 48 307
rect 48 306 49 307
rect 49 306 50 307
rect 50 306 51 307
rect 51 306 52 307
rect 52 306 53 307
rect 53 306 54 307
rect 54 306 55 307
rect 55 306 56 307
rect 105 306 106 307
rect 106 306 107 307
rect 107 306 108 307
rect 108 306 109 307
rect 109 306 110 307
rect 110 306 111 307
rect 111 306 112 307
rect 527 306 528 307
rect 528 306 529 307
rect 529 306 530 307
rect 530 306 531 307
rect 531 306 532 307
rect 532 306 533 307
rect 533 306 534 307
rect 534 306 535 307
rect 535 306 536 307
rect 536 306 537 307
rect 537 306 538 307
rect 538 306 539 307
rect 34 305 35 306
rect 35 305 36 306
rect 36 305 37 306
rect 37 305 38 306
rect 38 305 39 306
rect 39 305 40 306
rect 40 305 41 306
rect 41 305 42 306
rect 42 305 43 306
rect 43 305 44 306
rect 44 305 45 306
rect 45 305 46 306
rect 46 305 47 306
rect 47 305 48 306
rect 48 305 49 306
rect 49 305 50 306
rect 50 305 51 306
rect 51 305 52 306
rect 52 305 53 306
rect 53 305 54 306
rect 54 305 55 306
rect 55 305 56 306
rect 56 305 57 306
rect 57 305 58 306
rect 103 305 104 306
rect 104 305 105 306
rect 105 305 106 306
rect 106 305 107 306
rect 107 305 108 306
rect 108 305 109 306
rect 109 305 110 306
rect 110 305 111 306
rect 111 305 112 306
rect 527 305 528 306
rect 528 305 529 306
rect 529 305 530 306
rect 530 305 531 306
rect 531 305 532 306
rect 532 305 533 306
rect 533 305 534 306
rect 534 305 535 306
rect 535 305 536 306
rect 536 305 537 306
rect 537 305 538 306
rect 538 305 539 306
rect 34 304 35 305
rect 35 304 36 305
rect 36 304 37 305
rect 37 304 38 305
rect 38 304 39 305
rect 39 304 40 305
rect 40 304 41 305
rect 41 304 42 305
rect 42 304 43 305
rect 43 304 44 305
rect 44 304 45 305
rect 45 304 46 305
rect 46 304 47 305
rect 47 304 48 305
rect 48 304 49 305
rect 49 304 50 305
rect 50 304 51 305
rect 51 304 52 305
rect 52 304 53 305
rect 53 304 54 305
rect 54 304 55 305
rect 55 304 56 305
rect 56 304 57 305
rect 57 304 58 305
rect 103 304 104 305
rect 104 304 105 305
rect 105 304 106 305
rect 106 304 107 305
rect 107 304 108 305
rect 108 304 109 305
rect 109 304 110 305
rect 110 304 111 305
rect 111 304 112 305
rect 527 304 528 305
rect 528 304 529 305
rect 529 304 530 305
rect 530 304 531 305
rect 531 304 532 305
rect 532 304 533 305
rect 533 304 534 305
rect 534 304 535 305
rect 535 304 536 305
rect 536 304 537 305
rect 537 304 538 305
rect 538 304 539 305
rect 34 303 35 304
rect 35 303 36 304
rect 36 303 37 304
rect 37 303 38 304
rect 38 303 39 304
rect 39 303 40 304
rect 40 303 41 304
rect 41 303 42 304
rect 42 303 43 304
rect 43 303 44 304
rect 44 303 45 304
rect 45 303 46 304
rect 46 303 47 304
rect 47 303 48 304
rect 48 303 49 304
rect 49 303 50 304
rect 50 303 51 304
rect 51 303 52 304
rect 52 303 53 304
rect 53 303 54 304
rect 54 303 55 304
rect 55 303 56 304
rect 56 303 57 304
rect 57 303 58 304
rect 58 303 59 304
rect 103 303 104 304
rect 104 303 105 304
rect 105 303 106 304
rect 106 303 107 304
rect 107 303 108 304
rect 108 303 109 304
rect 109 303 110 304
rect 110 303 111 304
rect 111 303 112 304
rect 527 303 528 304
rect 528 303 529 304
rect 529 303 530 304
rect 530 303 531 304
rect 531 303 532 304
rect 532 303 533 304
rect 533 303 534 304
rect 534 303 535 304
rect 535 303 536 304
rect 536 303 537 304
rect 537 303 538 304
rect 538 303 539 304
rect 38 302 39 303
rect 39 302 40 303
rect 40 302 41 303
rect 41 302 42 303
rect 42 302 43 303
rect 43 302 44 303
rect 44 302 45 303
rect 45 302 46 303
rect 46 302 47 303
rect 47 302 48 303
rect 48 302 49 303
rect 49 302 50 303
rect 50 302 51 303
rect 51 302 52 303
rect 52 302 53 303
rect 53 302 54 303
rect 54 302 55 303
rect 55 302 56 303
rect 56 302 57 303
rect 57 302 58 303
rect 58 302 59 303
rect 103 302 104 303
rect 104 302 105 303
rect 105 302 106 303
rect 106 302 107 303
rect 107 302 108 303
rect 108 302 109 303
rect 109 302 110 303
rect 529 302 530 303
rect 530 302 531 303
rect 531 302 532 303
rect 532 302 533 303
rect 533 302 534 303
rect 534 302 535 303
rect 535 302 536 303
rect 536 302 537 303
rect 537 302 538 303
rect 538 302 539 303
rect 38 301 39 302
rect 39 301 40 302
rect 40 301 41 302
rect 41 301 42 302
rect 42 301 43 302
rect 43 301 44 302
rect 44 301 45 302
rect 45 301 46 302
rect 46 301 47 302
rect 47 301 48 302
rect 48 301 49 302
rect 49 301 50 302
rect 50 301 51 302
rect 51 301 52 302
rect 52 301 53 302
rect 53 301 54 302
rect 54 301 55 302
rect 55 301 56 302
rect 56 301 57 302
rect 57 301 58 302
rect 58 301 59 302
rect 59 301 60 302
rect 60 301 61 302
rect 61 301 62 302
rect 62 301 63 302
rect 102 301 103 302
rect 103 301 104 302
rect 104 301 105 302
rect 105 301 106 302
rect 106 301 107 302
rect 107 301 108 302
rect 108 301 109 302
rect 109 301 110 302
rect 118 301 119 302
rect 119 301 120 302
rect 120 301 121 302
rect 121 301 122 302
rect 122 301 123 302
rect 123 301 124 302
rect 124 301 125 302
rect 125 301 126 302
rect 126 301 127 302
rect 127 301 128 302
rect 128 301 129 302
rect 129 301 130 302
rect 130 301 131 302
rect 131 301 132 302
rect 132 301 133 302
rect 133 301 134 302
rect 134 301 135 302
rect 135 301 136 302
rect 136 301 137 302
rect 137 301 138 302
rect 138 301 139 302
rect 139 301 140 302
rect 140 301 141 302
rect 141 301 142 302
rect 142 301 143 302
rect 143 301 144 302
rect 144 301 145 302
rect 145 301 146 302
rect 150 301 151 302
rect 151 301 152 302
rect 152 301 153 302
rect 153 301 154 302
rect 154 301 155 302
rect 155 301 156 302
rect 156 301 157 302
rect 157 301 158 302
rect 158 301 159 302
rect 159 301 160 302
rect 160 301 161 302
rect 161 301 162 302
rect 162 301 163 302
rect 163 301 164 302
rect 164 301 165 302
rect 165 301 166 302
rect 166 301 167 302
rect 167 301 168 302
rect 168 301 169 302
rect 169 301 170 302
rect 170 301 171 302
rect 171 301 172 302
rect 172 301 173 302
rect 173 301 174 302
rect 174 301 175 302
rect 175 301 176 302
rect 176 301 177 302
rect 529 301 530 302
rect 530 301 531 302
rect 531 301 532 302
rect 532 301 533 302
rect 533 301 534 302
rect 534 301 535 302
rect 535 301 536 302
rect 536 301 537 302
rect 537 301 538 302
rect 538 301 539 302
rect 42 300 43 301
rect 43 300 44 301
rect 44 300 45 301
rect 45 300 46 301
rect 46 300 47 301
rect 47 300 48 301
rect 48 300 49 301
rect 49 300 50 301
rect 50 300 51 301
rect 51 300 52 301
rect 52 300 53 301
rect 53 300 54 301
rect 54 300 55 301
rect 55 300 56 301
rect 56 300 57 301
rect 57 300 58 301
rect 58 300 59 301
rect 59 300 60 301
rect 60 300 61 301
rect 61 300 62 301
rect 62 300 63 301
rect 102 300 103 301
rect 103 300 104 301
rect 104 300 105 301
rect 105 300 106 301
rect 106 300 107 301
rect 107 300 108 301
rect 108 300 109 301
rect 109 300 110 301
rect 118 300 119 301
rect 119 300 120 301
rect 120 300 121 301
rect 121 300 122 301
rect 122 300 123 301
rect 123 300 124 301
rect 124 300 125 301
rect 125 300 126 301
rect 126 300 127 301
rect 127 300 128 301
rect 128 300 129 301
rect 129 300 130 301
rect 130 300 131 301
rect 131 300 132 301
rect 132 300 133 301
rect 133 300 134 301
rect 134 300 135 301
rect 135 300 136 301
rect 136 300 137 301
rect 137 300 138 301
rect 138 300 139 301
rect 139 300 140 301
rect 140 300 141 301
rect 141 300 142 301
rect 142 300 143 301
rect 143 300 144 301
rect 144 300 145 301
rect 145 300 146 301
rect 150 300 151 301
rect 151 300 152 301
rect 152 300 153 301
rect 153 300 154 301
rect 154 300 155 301
rect 155 300 156 301
rect 156 300 157 301
rect 157 300 158 301
rect 158 300 159 301
rect 159 300 160 301
rect 160 300 161 301
rect 161 300 162 301
rect 162 300 163 301
rect 163 300 164 301
rect 164 300 165 301
rect 165 300 166 301
rect 166 300 167 301
rect 167 300 168 301
rect 168 300 169 301
rect 169 300 170 301
rect 170 300 171 301
rect 171 300 172 301
rect 172 300 173 301
rect 173 300 174 301
rect 174 300 175 301
rect 175 300 176 301
rect 176 300 177 301
rect 529 300 530 301
rect 530 300 531 301
rect 531 300 532 301
rect 532 300 533 301
rect 533 300 534 301
rect 534 300 535 301
rect 535 300 536 301
rect 536 300 537 301
rect 537 300 538 301
rect 538 300 539 301
rect 42 299 43 300
rect 43 299 44 300
rect 44 299 45 300
rect 45 299 46 300
rect 46 299 47 300
rect 47 299 48 300
rect 48 299 49 300
rect 49 299 50 300
rect 50 299 51 300
rect 51 299 52 300
rect 52 299 53 300
rect 53 299 54 300
rect 54 299 55 300
rect 55 299 56 300
rect 56 299 57 300
rect 57 299 58 300
rect 58 299 59 300
rect 59 299 60 300
rect 60 299 61 300
rect 61 299 62 300
rect 62 299 63 300
rect 63 299 64 300
rect 64 299 65 300
rect 100 299 101 300
rect 101 299 102 300
rect 102 299 103 300
rect 103 299 104 300
rect 104 299 105 300
rect 105 299 106 300
rect 106 299 107 300
rect 107 299 108 300
rect 108 299 109 300
rect 109 299 110 300
rect 118 299 119 300
rect 119 299 120 300
rect 120 299 121 300
rect 121 299 122 300
rect 122 299 123 300
rect 123 299 124 300
rect 124 299 125 300
rect 125 299 126 300
rect 126 299 127 300
rect 127 299 128 300
rect 128 299 129 300
rect 129 299 130 300
rect 130 299 131 300
rect 131 299 132 300
rect 132 299 133 300
rect 133 299 134 300
rect 134 299 135 300
rect 135 299 136 300
rect 136 299 137 300
rect 137 299 138 300
rect 138 299 139 300
rect 139 299 140 300
rect 140 299 141 300
rect 141 299 142 300
rect 142 299 143 300
rect 143 299 144 300
rect 144 299 145 300
rect 145 299 146 300
rect 150 299 151 300
rect 151 299 152 300
rect 152 299 153 300
rect 153 299 154 300
rect 154 299 155 300
rect 155 299 156 300
rect 156 299 157 300
rect 157 299 158 300
rect 158 299 159 300
rect 159 299 160 300
rect 160 299 161 300
rect 161 299 162 300
rect 162 299 163 300
rect 163 299 164 300
rect 164 299 165 300
rect 165 299 166 300
rect 166 299 167 300
rect 167 299 168 300
rect 168 299 169 300
rect 169 299 170 300
rect 170 299 171 300
rect 171 299 172 300
rect 172 299 173 300
rect 173 299 174 300
rect 174 299 175 300
rect 175 299 176 300
rect 176 299 177 300
rect 529 299 530 300
rect 530 299 531 300
rect 531 299 532 300
rect 532 299 533 300
rect 533 299 534 300
rect 534 299 535 300
rect 535 299 536 300
rect 536 299 537 300
rect 537 299 538 300
rect 538 299 539 300
rect 45 298 46 299
rect 46 298 47 299
rect 47 298 48 299
rect 48 298 49 299
rect 49 298 50 299
rect 50 298 51 299
rect 51 298 52 299
rect 52 298 53 299
rect 53 298 54 299
rect 54 298 55 299
rect 55 298 56 299
rect 56 298 57 299
rect 57 298 58 299
rect 58 298 59 299
rect 59 298 60 299
rect 60 298 61 299
rect 61 298 62 299
rect 62 298 63 299
rect 63 298 64 299
rect 64 298 65 299
rect 100 298 101 299
rect 101 298 102 299
rect 102 298 103 299
rect 103 298 104 299
rect 104 298 105 299
rect 105 298 106 299
rect 106 298 107 299
rect 107 298 108 299
rect 122 298 123 299
rect 123 298 124 299
rect 124 298 125 299
rect 125 298 126 299
rect 126 298 127 299
rect 127 298 128 299
rect 128 298 129 299
rect 129 298 130 299
rect 130 298 131 299
rect 131 298 132 299
rect 132 298 133 299
rect 133 298 134 299
rect 134 298 135 299
rect 135 298 136 299
rect 136 298 137 299
rect 137 298 138 299
rect 138 298 139 299
rect 139 298 140 299
rect 140 298 141 299
rect 141 298 142 299
rect 156 298 157 299
rect 157 298 158 299
rect 158 298 159 299
rect 159 298 160 299
rect 160 298 161 299
rect 161 298 162 299
rect 162 298 163 299
rect 163 298 164 299
rect 164 298 165 299
rect 165 298 166 299
rect 166 298 167 299
rect 167 298 168 299
rect 168 298 169 299
rect 169 298 170 299
rect 170 298 171 299
rect 171 298 172 299
rect 529 298 530 299
rect 530 298 531 299
rect 531 298 532 299
rect 532 298 533 299
rect 533 298 534 299
rect 534 298 535 299
rect 535 298 536 299
rect 536 298 537 299
rect 537 298 538 299
rect 538 298 539 299
rect 45 297 46 298
rect 46 297 47 298
rect 47 297 48 298
rect 48 297 49 298
rect 49 297 50 298
rect 50 297 51 298
rect 51 297 52 298
rect 52 297 53 298
rect 53 297 54 298
rect 54 297 55 298
rect 55 297 56 298
rect 56 297 57 298
rect 57 297 58 298
rect 58 297 59 298
rect 59 297 60 298
rect 60 297 61 298
rect 61 297 62 298
rect 62 297 63 298
rect 63 297 64 298
rect 64 297 65 298
rect 65 297 66 298
rect 66 297 67 298
rect 67 297 68 298
rect 68 297 69 298
rect 69 297 70 298
rect 70 297 71 298
rect 98 297 99 298
rect 99 297 100 298
rect 100 297 101 298
rect 101 297 102 298
rect 102 297 103 298
rect 103 297 104 298
rect 104 297 105 298
rect 105 297 106 298
rect 106 297 107 298
rect 107 297 108 298
rect 122 297 123 298
rect 123 297 124 298
rect 124 297 125 298
rect 125 297 126 298
rect 126 297 127 298
rect 127 297 128 298
rect 128 297 129 298
rect 129 297 130 298
rect 130 297 131 298
rect 131 297 132 298
rect 132 297 133 298
rect 133 297 134 298
rect 134 297 135 298
rect 135 297 136 298
rect 136 297 137 298
rect 137 297 138 298
rect 138 297 139 298
rect 139 297 140 298
rect 140 297 141 298
rect 141 297 142 298
rect 156 297 157 298
rect 157 297 158 298
rect 158 297 159 298
rect 159 297 160 298
rect 160 297 161 298
rect 161 297 162 298
rect 162 297 163 298
rect 163 297 164 298
rect 164 297 165 298
rect 165 297 166 298
rect 166 297 167 298
rect 167 297 168 298
rect 168 297 169 298
rect 169 297 170 298
rect 170 297 171 298
rect 171 297 172 298
rect 529 297 530 298
rect 530 297 531 298
rect 531 297 532 298
rect 532 297 533 298
rect 533 297 534 298
rect 534 297 535 298
rect 535 297 536 298
rect 536 297 537 298
rect 537 297 538 298
rect 538 297 539 298
rect 49 296 50 297
rect 50 296 51 297
rect 51 296 52 297
rect 52 296 53 297
rect 53 296 54 297
rect 54 296 55 297
rect 55 296 56 297
rect 56 296 57 297
rect 57 296 58 297
rect 58 296 59 297
rect 59 296 60 297
rect 60 296 61 297
rect 61 296 62 297
rect 62 296 63 297
rect 63 296 64 297
rect 64 296 65 297
rect 65 296 66 297
rect 66 296 67 297
rect 67 296 68 297
rect 68 296 69 297
rect 69 296 70 297
rect 70 296 71 297
rect 98 296 99 297
rect 99 296 100 297
rect 100 296 101 297
rect 101 296 102 297
rect 102 296 103 297
rect 103 296 104 297
rect 104 296 105 297
rect 105 296 106 297
rect 126 296 127 297
rect 127 296 128 297
rect 128 296 129 297
rect 129 296 130 297
rect 130 296 131 297
rect 131 296 132 297
rect 132 296 133 297
rect 133 296 134 297
rect 134 296 135 297
rect 135 296 136 297
rect 136 296 137 297
rect 137 296 138 297
rect 160 296 161 297
rect 161 296 162 297
rect 162 296 163 297
rect 163 296 164 297
rect 164 296 165 297
rect 165 296 166 297
rect 166 296 167 297
rect 167 296 168 297
rect 168 296 169 297
rect 169 296 170 297
rect 529 296 530 297
rect 530 296 531 297
rect 531 296 532 297
rect 532 296 533 297
rect 533 296 534 297
rect 534 296 535 297
rect 535 296 536 297
rect 536 296 537 297
rect 537 296 538 297
rect 538 296 539 297
rect 49 295 50 296
rect 50 295 51 296
rect 51 295 52 296
rect 52 295 53 296
rect 53 295 54 296
rect 54 295 55 296
rect 55 295 56 296
rect 56 295 57 296
rect 57 295 58 296
rect 58 295 59 296
rect 59 295 60 296
rect 60 295 61 296
rect 61 295 62 296
rect 62 295 63 296
rect 63 295 64 296
rect 64 295 65 296
rect 65 295 66 296
rect 66 295 67 296
rect 67 295 68 296
rect 68 295 69 296
rect 69 295 70 296
rect 70 295 71 296
rect 71 295 72 296
rect 72 295 73 296
rect 73 295 74 296
rect 96 295 97 296
rect 97 295 98 296
rect 98 295 99 296
rect 99 295 100 296
rect 100 295 101 296
rect 101 295 102 296
rect 102 295 103 296
rect 103 295 104 296
rect 104 295 105 296
rect 105 295 106 296
rect 126 295 127 296
rect 127 295 128 296
rect 128 295 129 296
rect 129 295 130 296
rect 130 295 131 296
rect 131 295 132 296
rect 132 295 133 296
rect 133 295 134 296
rect 134 295 135 296
rect 135 295 136 296
rect 136 295 137 296
rect 137 295 138 296
rect 158 295 159 296
rect 159 295 160 296
rect 160 295 161 296
rect 161 295 162 296
rect 162 295 163 296
rect 163 295 164 296
rect 164 295 165 296
rect 165 295 166 296
rect 166 295 167 296
rect 167 295 168 296
rect 168 295 169 296
rect 169 295 170 296
rect 529 295 530 296
rect 530 295 531 296
rect 531 295 532 296
rect 532 295 533 296
rect 533 295 534 296
rect 534 295 535 296
rect 535 295 536 296
rect 536 295 537 296
rect 537 295 538 296
rect 538 295 539 296
rect 53 294 54 295
rect 54 294 55 295
rect 55 294 56 295
rect 56 294 57 295
rect 57 294 58 295
rect 58 294 59 295
rect 59 294 60 295
rect 60 294 61 295
rect 61 294 62 295
rect 62 294 63 295
rect 63 294 64 295
rect 64 294 65 295
rect 65 294 66 295
rect 66 294 67 295
rect 67 294 68 295
rect 68 294 69 295
rect 69 294 70 295
rect 70 294 71 295
rect 71 294 72 295
rect 72 294 73 295
rect 73 294 74 295
rect 96 294 97 295
rect 97 294 98 295
rect 98 294 99 295
rect 99 294 100 295
rect 100 294 101 295
rect 101 294 102 295
rect 102 294 103 295
rect 103 294 104 295
rect 104 294 105 295
rect 105 294 106 295
rect 126 294 127 295
rect 127 294 128 295
rect 128 294 129 295
rect 129 294 130 295
rect 130 294 131 295
rect 131 294 132 295
rect 132 294 133 295
rect 133 294 134 295
rect 134 294 135 295
rect 135 294 136 295
rect 136 294 137 295
rect 137 294 138 295
rect 158 294 159 295
rect 159 294 160 295
rect 160 294 161 295
rect 161 294 162 295
rect 162 294 163 295
rect 163 294 164 295
rect 164 294 165 295
rect 165 294 166 295
rect 529 294 530 295
rect 530 294 531 295
rect 531 294 532 295
rect 532 294 533 295
rect 533 294 534 295
rect 534 294 535 295
rect 535 294 536 295
rect 536 294 537 295
rect 537 294 538 295
rect 538 294 539 295
rect 53 293 54 294
rect 54 293 55 294
rect 55 293 56 294
rect 56 293 57 294
rect 57 293 58 294
rect 58 293 59 294
rect 59 293 60 294
rect 60 293 61 294
rect 61 293 62 294
rect 62 293 63 294
rect 63 293 64 294
rect 64 293 65 294
rect 65 293 66 294
rect 66 293 67 294
rect 67 293 68 294
rect 68 293 69 294
rect 69 293 70 294
rect 70 293 71 294
rect 71 293 72 294
rect 72 293 73 294
rect 73 293 74 294
rect 74 293 75 294
rect 75 293 76 294
rect 76 293 77 294
rect 77 293 78 294
rect 78 293 79 294
rect 79 293 80 294
rect 80 293 81 294
rect 81 293 82 294
rect 82 293 83 294
rect 83 293 84 294
rect 92 293 93 294
rect 93 293 94 294
rect 94 293 95 294
rect 95 293 96 294
rect 96 293 97 294
rect 97 293 98 294
rect 98 293 99 294
rect 99 293 100 294
rect 100 293 101 294
rect 101 293 102 294
rect 102 293 103 294
rect 103 293 104 294
rect 104 293 105 294
rect 105 293 106 294
rect 126 293 127 294
rect 127 293 128 294
rect 128 293 129 294
rect 129 293 130 294
rect 130 293 131 294
rect 131 293 132 294
rect 132 293 133 294
rect 133 293 134 294
rect 134 293 135 294
rect 135 293 136 294
rect 136 293 137 294
rect 137 293 138 294
rect 158 293 159 294
rect 159 293 160 294
rect 160 293 161 294
rect 161 293 162 294
rect 162 293 163 294
rect 163 293 164 294
rect 164 293 165 294
rect 165 293 166 294
rect 529 293 530 294
rect 530 293 531 294
rect 531 293 532 294
rect 532 293 533 294
rect 533 293 534 294
rect 534 293 535 294
rect 535 293 536 294
rect 536 293 537 294
rect 537 293 538 294
rect 538 293 539 294
rect 57 292 58 293
rect 58 292 59 293
rect 59 292 60 293
rect 60 292 61 293
rect 61 292 62 293
rect 62 292 63 293
rect 63 292 64 293
rect 64 292 65 293
rect 65 292 66 293
rect 66 292 67 293
rect 67 292 68 293
rect 68 292 69 293
rect 69 292 70 293
rect 70 292 71 293
rect 71 292 72 293
rect 72 292 73 293
rect 73 292 74 293
rect 74 292 75 293
rect 75 292 76 293
rect 76 292 77 293
rect 77 292 78 293
rect 78 292 79 293
rect 79 292 80 293
rect 80 292 81 293
rect 81 292 82 293
rect 82 292 83 293
rect 83 292 84 293
rect 92 292 93 293
rect 93 292 94 293
rect 94 292 95 293
rect 95 292 96 293
rect 96 292 97 293
rect 97 292 98 293
rect 98 292 99 293
rect 99 292 100 293
rect 100 292 101 293
rect 101 292 102 293
rect 102 292 103 293
rect 103 292 104 293
rect 126 292 127 293
rect 127 292 128 293
rect 128 292 129 293
rect 129 292 130 293
rect 130 292 131 293
rect 131 292 132 293
rect 132 292 133 293
rect 133 292 134 293
rect 134 292 135 293
rect 135 292 136 293
rect 136 292 137 293
rect 137 292 138 293
rect 158 292 159 293
rect 159 292 160 293
rect 160 292 161 293
rect 161 292 162 293
rect 162 292 163 293
rect 163 292 164 293
rect 530 292 531 293
rect 531 292 532 293
rect 532 292 533 293
rect 533 292 534 293
rect 534 292 535 293
rect 535 292 536 293
rect 536 292 537 293
rect 537 292 538 293
rect 538 292 539 293
rect 57 291 58 292
rect 58 291 59 292
rect 59 291 60 292
rect 60 291 61 292
rect 61 291 62 292
rect 62 291 63 292
rect 63 291 64 292
rect 64 291 65 292
rect 65 291 66 292
rect 66 291 67 292
rect 67 291 68 292
rect 68 291 69 292
rect 69 291 70 292
rect 70 291 71 292
rect 71 291 72 292
rect 72 291 73 292
rect 73 291 74 292
rect 74 291 75 292
rect 75 291 76 292
rect 76 291 77 292
rect 77 291 78 292
rect 78 291 79 292
rect 79 291 80 292
rect 80 291 81 292
rect 81 291 82 292
rect 82 291 83 292
rect 83 291 84 292
rect 84 291 85 292
rect 85 291 86 292
rect 86 291 87 292
rect 87 291 88 292
rect 88 291 89 292
rect 89 291 90 292
rect 90 291 91 292
rect 91 291 92 292
rect 92 291 93 292
rect 93 291 94 292
rect 94 291 95 292
rect 95 291 96 292
rect 96 291 97 292
rect 97 291 98 292
rect 98 291 99 292
rect 99 291 100 292
rect 100 291 101 292
rect 101 291 102 292
rect 102 291 103 292
rect 103 291 104 292
rect 126 291 127 292
rect 127 291 128 292
rect 128 291 129 292
rect 129 291 130 292
rect 130 291 131 292
rect 131 291 132 292
rect 132 291 133 292
rect 133 291 134 292
rect 134 291 135 292
rect 135 291 136 292
rect 136 291 137 292
rect 137 291 138 292
rect 156 291 157 292
rect 157 291 158 292
rect 158 291 159 292
rect 159 291 160 292
rect 160 291 161 292
rect 161 291 162 292
rect 162 291 163 292
rect 163 291 164 292
rect 530 291 531 292
rect 531 291 532 292
rect 532 291 533 292
rect 533 291 534 292
rect 534 291 535 292
rect 535 291 536 292
rect 536 291 537 292
rect 537 291 538 292
rect 538 291 539 292
rect 62 290 63 291
rect 63 290 64 291
rect 64 290 65 291
rect 65 290 66 291
rect 66 290 67 291
rect 67 290 68 291
rect 68 290 69 291
rect 69 290 70 291
rect 70 290 71 291
rect 71 290 72 291
rect 72 290 73 291
rect 73 290 74 291
rect 74 290 75 291
rect 75 290 76 291
rect 76 290 77 291
rect 77 290 78 291
rect 78 290 79 291
rect 79 290 80 291
rect 80 290 81 291
rect 81 290 82 291
rect 82 290 83 291
rect 83 290 84 291
rect 84 290 85 291
rect 85 290 86 291
rect 86 290 87 291
rect 87 290 88 291
rect 88 290 89 291
rect 89 290 90 291
rect 90 290 91 291
rect 91 290 92 291
rect 92 290 93 291
rect 93 290 94 291
rect 94 290 95 291
rect 95 290 96 291
rect 96 290 97 291
rect 97 290 98 291
rect 98 290 99 291
rect 99 290 100 291
rect 100 290 101 291
rect 101 290 102 291
rect 102 290 103 291
rect 103 290 104 291
rect 126 290 127 291
rect 127 290 128 291
rect 128 290 129 291
rect 129 290 130 291
rect 130 290 131 291
rect 131 290 132 291
rect 132 290 133 291
rect 133 290 134 291
rect 134 290 135 291
rect 135 290 136 291
rect 156 290 157 291
rect 157 290 158 291
rect 158 290 159 291
rect 159 290 160 291
rect 160 290 161 291
rect 161 290 162 291
rect 162 290 163 291
rect 530 290 531 291
rect 531 290 532 291
rect 532 290 533 291
rect 533 290 534 291
rect 534 290 535 291
rect 535 290 536 291
rect 536 290 537 291
rect 537 290 538 291
rect 538 290 539 291
rect 62 289 63 290
rect 63 289 64 290
rect 64 289 65 290
rect 65 289 66 290
rect 66 289 67 290
rect 67 289 68 290
rect 68 289 69 290
rect 69 289 70 290
rect 70 289 71 290
rect 71 289 72 290
rect 72 289 73 290
rect 73 289 74 290
rect 74 289 75 290
rect 75 289 76 290
rect 76 289 77 290
rect 77 289 78 290
rect 78 289 79 290
rect 79 289 80 290
rect 80 289 81 290
rect 81 289 82 290
rect 82 289 83 290
rect 83 289 84 290
rect 84 289 85 290
rect 85 289 86 290
rect 86 289 87 290
rect 87 289 88 290
rect 88 289 89 290
rect 89 289 90 290
rect 90 289 91 290
rect 91 289 92 290
rect 92 289 93 290
rect 93 289 94 290
rect 94 289 95 290
rect 95 289 96 290
rect 96 289 97 290
rect 97 289 98 290
rect 98 289 99 290
rect 99 289 100 290
rect 100 289 101 290
rect 101 289 102 290
rect 102 289 103 290
rect 103 289 104 290
rect 126 289 127 290
rect 127 289 128 290
rect 128 289 129 290
rect 129 289 130 290
rect 130 289 131 290
rect 131 289 132 290
rect 132 289 133 290
rect 133 289 134 290
rect 134 289 135 290
rect 135 289 136 290
rect 154 289 155 290
rect 155 289 156 290
rect 156 289 157 290
rect 157 289 158 290
rect 158 289 159 290
rect 159 289 160 290
rect 160 289 161 290
rect 161 289 162 290
rect 162 289 163 290
rect 530 289 531 290
rect 531 289 532 290
rect 532 289 533 290
rect 533 289 534 290
rect 534 289 535 290
rect 535 289 536 290
rect 536 289 537 290
rect 537 289 538 290
rect 538 289 539 290
rect 66 288 67 289
rect 67 288 68 289
rect 68 288 69 289
rect 69 288 70 289
rect 70 288 71 289
rect 71 288 72 289
rect 72 288 73 289
rect 73 288 74 289
rect 74 288 75 289
rect 75 288 76 289
rect 76 288 77 289
rect 77 288 78 289
rect 78 288 79 289
rect 79 288 80 289
rect 80 288 81 289
rect 81 288 82 289
rect 82 288 83 289
rect 83 288 84 289
rect 84 288 85 289
rect 85 288 86 289
rect 86 288 87 289
rect 87 288 88 289
rect 88 288 89 289
rect 89 288 90 289
rect 90 288 91 289
rect 91 288 92 289
rect 92 288 93 289
rect 93 288 94 289
rect 94 288 95 289
rect 95 288 96 289
rect 96 288 97 289
rect 97 288 98 289
rect 98 288 99 289
rect 99 288 100 289
rect 100 288 101 289
rect 101 288 102 289
rect 102 288 103 289
rect 103 288 104 289
rect 126 288 127 289
rect 127 288 128 289
rect 128 288 129 289
rect 129 288 130 289
rect 130 288 131 289
rect 131 288 132 289
rect 132 288 133 289
rect 133 288 134 289
rect 134 288 135 289
rect 135 288 136 289
rect 154 288 155 289
rect 155 288 156 289
rect 156 288 157 289
rect 157 288 158 289
rect 158 288 159 289
rect 159 288 160 289
rect 160 288 161 289
rect 530 288 531 289
rect 531 288 532 289
rect 532 288 533 289
rect 533 288 534 289
rect 534 288 535 289
rect 535 288 536 289
rect 536 288 537 289
rect 537 288 538 289
rect 538 288 539 289
rect 66 287 67 288
rect 67 287 68 288
rect 68 287 69 288
rect 69 287 70 288
rect 70 287 71 288
rect 71 287 72 288
rect 72 287 73 288
rect 73 287 74 288
rect 74 287 75 288
rect 75 287 76 288
rect 76 287 77 288
rect 77 287 78 288
rect 78 287 79 288
rect 79 287 80 288
rect 80 287 81 288
rect 81 287 82 288
rect 82 287 83 288
rect 83 287 84 288
rect 84 287 85 288
rect 85 287 86 288
rect 86 287 87 288
rect 87 287 88 288
rect 88 287 89 288
rect 89 287 90 288
rect 90 287 91 288
rect 91 287 92 288
rect 92 287 93 288
rect 93 287 94 288
rect 94 287 95 288
rect 95 287 96 288
rect 96 287 97 288
rect 97 287 98 288
rect 98 287 99 288
rect 99 287 100 288
rect 100 287 101 288
rect 101 287 102 288
rect 102 287 103 288
rect 103 287 104 288
rect 126 287 127 288
rect 127 287 128 288
rect 128 287 129 288
rect 129 287 130 288
rect 130 287 131 288
rect 131 287 132 288
rect 132 287 133 288
rect 133 287 134 288
rect 134 287 135 288
rect 135 287 136 288
rect 136 287 137 288
rect 137 287 138 288
rect 152 287 153 288
rect 153 287 154 288
rect 154 287 155 288
rect 155 287 156 288
rect 156 287 157 288
rect 157 287 158 288
rect 158 287 159 288
rect 159 287 160 288
rect 160 287 161 288
rect 530 287 531 288
rect 531 287 532 288
rect 532 287 533 288
rect 533 287 534 288
rect 534 287 535 288
rect 535 287 536 288
rect 536 287 537 288
rect 537 287 538 288
rect 538 287 539 288
rect 70 286 71 287
rect 71 286 72 287
rect 72 286 73 287
rect 73 286 74 287
rect 74 286 75 287
rect 75 286 76 287
rect 76 286 77 287
rect 77 286 78 287
rect 78 286 79 287
rect 79 286 80 287
rect 80 286 81 287
rect 81 286 82 287
rect 82 286 83 287
rect 83 286 84 287
rect 84 286 85 287
rect 85 286 86 287
rect 86 286 87 287
rect 87 286 88 287
rect 88 286 89 287
rect 89 286 90 287
rect 90 286 91 287
rect 91 286 92 287
rect 92 286 93 287
rect 93 286 94 287
rect 94 286 95 287
rect 95 286 96 287
rect 96 286 97 287
rect 97 286 98 287
rect 98 286 99 287
rect 99 286 100 287
rect 100 286 101 287
rect 101 286 102 287
rect 102 286 103 287
rect 126 286 127 287
rect 127 286 128 287
rect 128 286 129 287
rect 129 286 130 287
rect 130 286 131 287
rect 131 286 132 287
rect 132 286 133 287
rect 133 286 134 287
rect 134 286 135 287
rect 135 286 136 287
rect 136 286 137 287
rect 137 286 138 287
rect 152 286 153 287
rect 153 286 154 287
rect 154 286 155 287
rect 155 286 156 287
rect 156 286 157 287
rect 157 286 158 287
rect 158 286 159 287
rect 530 286 531 287
rect 531 286 532 287
rect 532 286 533 287
rect 533 286 534 287
rect 534 286 535 287
rect 535 286 536 287
rect 536 286 537 287
rect 537 286 538 287
rect 538 286 539 287
rect 70 285 71 286
rect 71 285 72 286
rect 72 285 73 286
rect 73 285 74 286
rect 74 285 75 286
rect 75 285 76 286
rect 76 285 77 286
rect 77 285 78 286
rect 78 285 79 286
rect 79 285 80 286
rect 80 285 81 286
rect 81 285 82 286
rect 82 285 83 286
rect 83 285 84 286
rect 84 285 85 286
rect 85 285 86 286
rect 86 285 87 286
rect 87 285 88 286
rect 88 285 89 286
rect 89 285 90 286
rect 90 285 91 286
rect 91 285 92 286
rect 92 285 93 286
rect 93 285 94 286
rect 94 285 95 286
rect 95 285 96 286
rect 96 285 97 286
rect 97 285 98 286
rect 98 285 99 286
rect 99 285 100 286
rect 100 285 101 286
rect 101 285 102 286
rect 102 285 103 286
rect 126 285 127 286
rect 127 285 128 286
rect 128 285 129 286
rect 129 285 130 286
rect 130 285 131 286
rect 131 285 132 286
rect 132 285 133 286
rect 133 285 134 286
rect 134 285 135 286
rect 135 285 136 286
rect 136 285 137 286
rect 137 285 138 286
rect 148 285 149 286
rect 149 285 150 286
rect 150 285 151 286
rect 151 285 152 286
rect 152 285 153 286
rect 153 285 154 286
rect 154 285 155 286
rect 155 285 156 286
rect 156 285 157 286
rect 157 285 158 286
rect 158 285 159 286
rect 530 285 531 286
rect 531 285 532 286
rect 532 285 533 286
rect 533 285 534 286
rect 534 285 535 286
rect 535 285 536 286
rect 536 285 537 286
rect 537 285 538 286
rect 538 285 539 286
rect 73 284 74 285
rect 74 284 75 285
rect 75 284 76 285
rect 76 284 77 285
rect 77 284 78 285
rect 78 284 79 285
rect 79 284 80 285
rect 80 284 81 285
rect 81 284 82 285
rect 82 284 83 285
rect 83 284 84 285
rect 84 284 85 285
rect 85 284 86 285
rect 86 284 87 285
rect 87 284 88 285
rect 88 284 89 285
rect 89 284 90 285
rect 90 284 91 285
rect 91 284 92 285
rect 92 284 93 285
rect 93 284 94 285
rect 94 284 95 285
rect 95 284 96 285
rect 96 284 97 285
rect 97 284 98 285
rect 98 284 99 285
rect 99 284 100 285
rect 100 284 101 285
rect 101 284 102 285
rect 102 284 103 285
rect 126 284 127 285
rect 127 284 128 285
rect 128 284 129 285
rect 129 284 130 285
rect 130 284 131 285
rect 131 284 132 285
rect 132 284 133 285
rect 133 284 134 285
rect 134 284 135 285
rect 135 284 136 285
rect 136 284 137 285
rect 137 284 138 285
rect 148 284 149 285
rect 149 284 150 285
rect 150 284 151 285
rect 151 284 152 285
rect 152 284 153 285
rect 153 284 154 285
rect 154 284 155 285
rect 155 284 156 285
rect 156 284 157 285
rect 530 284 531 285
rect 531 284 532 285
rect 532 284 533 285
rect 533 284 534 285
rect 534 284 535 285
rect 535 284 536 285
rect 536 284 537 285
rect 537 284 538 285
rect 538 284 539 285
rect 73 283 74 284
rect 74 283 75 284
rect 75 283 76 284
rect 76 283 77 284
rect 77 283 78 284
rect 78 283 79 284
rect 79 283 80 284
rect 80 283 81 284
rect 81 283 82 284
rect 82 283 83 284
rect 83 283 84 284
rect 84 283 85 284
rect 85 283 86 284
rect 86 283 87 284
rect 87 283 88 284
rect 88 283 89 284
rect 89 283 90 284
rect 90 283 91 284
rect 91 283 92 284
rect 92 283 93 284
rect 93 283 94 284
rect 94 283 95 284
rect 95 283 96 284
rect 96 283 97 284
rect 97 283 98 284
rect 98 283 99 284
rect 99 283 100 284
rect 100 283 101 284
rect 101 283 102 284
rect 102 283 103 284
rect 126 283 127 284
rect 127 283 128 284
rect 128 283 129 284
rect 129 283 130 284
rect 130 283 131 284
rect 131 283 132 284
rect 132 283 133 284
rect 133 283 134 284
rect 134 283 135 284
rect 135 283 136 284
rect 136 283 137 284
rect 137 283 138 284
rect 148 283 149 284
rect 149 283 150 284
rect 150 283 151 284
rect 151 283 152 284
rect 152 283 153 284
rect 153 283 154 284
rect 154 283 155 284
rect 155 283 156 284
rect 156 283 157 284
rect 530 283 531 284
rect 531 283 532 284
rect 532 283 533 284
rect 533 283 534 284
rect 534 283 535 284
rect 535 283 536 284
rect 536 283 537 284
rect 537 283 538 284
rect 538 283 539 284
rect 77 282 78 283
rect 78 282 79 283
rect 79 282 80 283
rect 80 282 81 283
rect 81 282 82 283
rect 82 282 83 283
rect 83 282 84 283
rect 84 282 85 283
rect 85 282 86 283
rect 86 282 87 283
rect 87 282 88 283
rect 88 282 89 283
rect 89 282 90 283
rect 90 282 91 283
rect 91 282 92 283
rect 92 282 93 283
rect 93 282 94 283
rect 94 282 95 283
rect 95 282 96 283
rect 96 282 97 283
rect 97 282 98 283
rect 98 282 99 283
rect 99 282 100 283
rect 100 282 101 283
rect 126 282 127 283
rect 127 282 128 283
rect 128 282 129 283
rect 129 282 130 283
rect 130 282 131 283
rect 131 282 132 283
rect 132 282 133 283
rect 133 282 134 283
rect 134 282 135 283
rect 135 282 136 283
rect 148 282 149 283
rect 149 282 150 283
rect 150 282 151 283
rect 151 282 152 283
rect 152 282 153 283
rect 153 282 154 283
rect 154 282 155 283
rect 530 282 531 283
rect 531 282 532 283
rect 532 282 533 283
rect 533 282 534 283
rect 534 282 535 283
rect 535 282 536 283
rect 536 282 537 283
rect 537 282 538 283
rect 538 282 539 283
rect 77 281 78 282
rect 78 281 79 282
rect 79 281 80 282
rect 80 281 81 282
rect 81 281 82 282
rect 82 281 83 282
rect 83 281 84 282
rect 84 281 85 282
rect 85 281 86 282
rect 86 281 87 282
rect 87 281 88 282
rect 88 281 89 282
rect 89 281 90 282
rect 90 281 91 282
rect 91 281 92 282
rect 92 281 93 282
rect 93 281 94 282
rect 94 281 95 282
rect 95 281 96 282
rect 96 281 97 282
rect 97 281 98 282
rect 98 281 99 282
rect 99 281 100 282
rect 100 281 101 282
rect 126 281 127 282
rect 127 281 128 282
rect 128 281 129 282
rect 129 281 130 282
rect 130 281 131 282
rect 131 281 132 282
rect 132 281 133 282
rect 133 281 134 282
rect 134 281 135 282
rect 135 281 136 282
rect 148 281 149 282
rect 149 281 150 282
rect 150 281 151 282
rect 151 281 152 282
rect 152 281 153 282
rect 153 281 154 282
rect 154 281 155 282
rect 530 281 531 282
rect 531 281 532 282
rect 532 281 533 282
rect 533 281 534 282
rect 534 281 535 282
rect 535 281 536 282
rect 536 281 537 282
rect 537 281 538 282
rect 538 281 539 282
rect 77 280 78 281
rect 78 280 79 281
rect 79 280 80 281
rect 80 280 81 281
rect 81 280 82 281
rect 82 280 83 281
rect 83 280 84 281
rect 84 280 85 281
rect 85 280 86 281
rect 86 280 87 281
rect 87 280 88 281
rect 88 280 89 281
rect 89 280 90 281
rect 90 280 91 281
rect 91 280 92 281
rect 92 280 93 281
rect 93 280 94 281
rect 94 280 95 281
rect 95 280 96 281
rect 96 280 97 281
rect 97 280 98 281
rect 98 280 99 281
rect 99 280 100 281
rect 100 280 101 281
rect 126 280 127 281
rect 127 280 128 281
rect 128 280 129 281
rect 129 280 130 281
rect 130 280 131 281
rect 131 280 132 281
rect 132 280 133 281
rect 133 280 134 281
rect 134 280 135 281
rect 135 280 136 281
rect 136 280 137 281
rect 137 280 138 281
rect 147 280 148 281
rect 148 280 149 281
rect 149 280 150 281
rect 150 280 151 281
rect 151 280 152 281
rect 152 280 153 281
rect 153 280 154 281
rect 154 280 155 281
rect 471 280 472 281
rect 472 280 473 281
rect 476 280 477 281
rect 477 280 478 281
rect 478 280 479 281
rect 480 280 481 281
rect 481 280 482 281
rect 482 280 483 281
rect 483 280 484 281
rect 484 280 485 281
rect 489 280 490 281
rect 490 280 491 281
rect 491 280 492 281
rect 530 280 531 281
rect 531 280 532 281
rect 532 280 533 281
rect 533 280 534 281
rect 534 280 535 281
rect 535 280 536 281
rect 536 280 537 281
rect 537 280 538 281
rect 538 280 539 281
rect 81 279 82 280
rect 82 279 83 280
rect 83 279 84 280
rect 84 279 85 280
rect 85 279 86 280
rect 86 279 87 280
rect 87 279 88 280
rect 88 279 89 280
rect 89 279 90 280
rect 90 279 91 280
rect 91 279 92 280
rect 92 279 93 280
rect 93 279 94 280
rect 94 279 95 280
rect 95 279 96 280
rect 96 279 97 280
rect 97 279 98 280
rect 98 279 99 280
rect 99 279 100 280
rect 100 279 101 280
rect 126 279 127 280
rect 127 279 128 280
rect 128 279 129 280
rect 129 279 130 280
rect 130 279 131 280
rect 131 279 132 280
rect 132 279 133 280
rect 133 279 134 280
rect 134 279 135 280
rect 135 279 136 280
rect 136 279 137 280
rect 137 279 138 280
rect 147 279 148 280
rect 148 279 149 280
rect 149 279 150 280
rect 150 279 151 280
rect 151 279 152 280
rect 152 279 153 280
rect 471 279 472 280
rect 472 279 473 280
rect 476 279 477 280
rect 477 279 478 280
rect 478 279 479 280
rect 480 279 481 280
rect 481 279 482 280
rect 482 279 483 280
rect 483 279 484 280
rect 484 279 485 280
rect 489 279 490 280
rect 490 279 491 280
rect 491 279 492 280
rect 532 279 533 280
rect 533 279 534 280
rect 534 279 535 280
rect 535 279 536 280
rect 536 279 537 280
rect 537 279 538 280
rect 538 279 539 280
rect 81 278 82 279
rect 82 278 83 279
rect 83 278 84 279
rect 84 278 85 279
rect 85 278 86 279
rect 86 278 87 279
rect 87 278 88 279
rect 88 278 89 279
rect 89 278 90 279
rect 90 278 91 279
rect 91 278 92 279
rect 92 278 93 279
rect 93 278 94 279
rect 94 278 95 279
rect 95 278 96 279
rect 96 278 97 279
rect 97 278 98 279
rect 98 278 99 279
rect 99 278 100 279
rect 100 278 101 279
rect 126 278 127 279
rect 127 278 128 279
rect 128 278 129 279
rect 129 278 130 279
rect 130 278 131 279
rect 131 278 132 279
rect 132 278 133 279
rect 133 278 134 279
rect 134 278 135 279
rect 135 278 136 279
rect 136 278 137 279
rect 137 278 138 279
rect 143 278 144 279
rect 144 278 145 279
rect 145 278 146 279
rect 146 278 147 279
rect 147 278 148 279
rect 148 278 149 279
rect 149 278 150 279
rect 150 278 151 279
rect 151 278 152 279
rect 152 278 153 279
rect 469 278 470 279
rect 470 278 471 279
rect 471 278 472 279
rect 472 278 473 279
rect 473 278 474 279
rect 474 278 475 279
rect 475 278 476 279
rect 476 278 477 279
rect 477 278 478 279
rect 478 278 479 279
rect 479 278 480 279
rect 480 278 481 279
rect 481 278 482 279
rect 482 278 483 279
rect 483 278 484 279
rect 484 278 485 279
rect 485 278 486 279
rect 486 278 487 279
rect 487 278 488 279
rect 488 278 489 279
rect 489 278 490 279
rect 490 278 491 279
rect 491 278 492 279
rect 492 278 493 279
rect 493 278 494 279
rect 494 278 495 279
rect 495 278 496 279
rect 530 278 531 279
rect 531 278 532 279
rect 532 278 533 279
rect 533 278 534 279
rect 534 278 535 279
rect 535 278 536 279
rect 536 278 537 279
rect 537 278 538 279
rect 538 278 539 279
rect 83 277 84 278
rect 84 277 85 278
rect 85 277 86 278
rect 86 277 87 278
rect 87 277 88 278
rect 88 277 89 278
rect 89 277 90 278
rect 90 277 91 278
rect 91 277 92 278
rect 92 277 93 278
rect 93 277 94 278
rect 94 277 95 278
rect 95 277 96 278
rect 96 277 97 278
rect 97 277 98 278
rect 98 277 99 278
rect 99 277 100 278
rect 100 277 101 278
rect 126 277 127 278
rect 127 277 128 278
rect 128 277 129 278
rect 129 277 130 278
rect 130 277 131 278
rect 131 277 132 278
rect 132 277 133 278
rect 133 277 134 278
rect 134 277 135 278
rect 135 277 136 278
rect 136 277 137 278
rect 137 277 138 278
rect 143 277 144 278
rect 144 277 145 278
rect 145 277 146 278
rect 146 277 147 278
rect 147 277 148 278
rect 148 277 149 278
rect 149 277 150 278
rect 150 277 151 278
rect 469 277 470 278
rect 470 277 471 278
rect 471 277 472 278
rect 472 277 473 278
rect 473 277 474 278
rect 474 277 475 278
rect 475 277 476 278
rect 476 277 477 278
rect 477 277 478 278
rect 478 277 479 278
rect 479 277 480 278
rect 480 277 481 278
rect 481 277 482 278
rect 482 277 483 278
rect 483 277 484 278
rect 484 277 485 278
rect 485 277 486 278
rect 486 277 487 278
rect 487 277 488 278
rect 488 277 489 278
rect 489 277 490 278
rect 490 277 491 278
rect 491 277 492 278
rect 492 277 493 278
rect 493 277 494 278
rect 494 277 495 278
rect 495 277 496 278
rect 530 277 531 278
rect 531 277 532 278
rect 532 277 533 278
rect 533 277 534 278
rect 534 277 535 278
rect 535 277 536 278
rect 536 277 537 278
rect 537 277 538 278
rect 538 277 539 278
rect 83 276 84 277
rect 84 276 85 277
rect 85 276 86 277
rect 86 276 87 277
rect 87 276 88 277
rect 88 276 89 277
rect 89 276 90 277
rect 90 276 91 277
rect 91 276 92 277
rect 92 276 93 277
rect 93 276 94 277
rect 94 276 95 277
rect 95 276 96 277
rect 96 276 97 277
rect 97 276 98 277
rect 98 276 99 277
rect 99 276 100 277
rect 100 276 101 277
rect 126 276 127 277
rect 127 276 128 277
rect 128 276 129 277
rect 129 276 130 277
rect 130 276 131 277
rect 131 276 132 277
rect 132 276 133 277
rect 133 276 134 277
rect 134 276 135 277
rect 135 276 136 277
rect 136 276 137 277
rect 137 276 138 277
rect 141 276 142 277
rect 142 276 143 277
rect 143 276 144 277
rect 144 276 145 277
rect 145 276 146 277
rect 146 276 147 277
rect 147 276 148 277
rect 148 276 149 277
rect 149 276 150 277
rect 150 276 151 277
rect 469 276 470 277
rect 470 276 471 277
rect 471 276 472 277
rect 472 276 473 277
rect 473 276 474 277
rect 474 276 475 277
rect 475 276 476 277
rect 476 276 477 277
rect 477 276 478 277
rect 478 276 479 277
rect 479 276 480 277
rect 480 276 481 277
rect 481 276 482 277
rect 482 276 483 277
rect 483 276 484 277
rect 484 276 485 277
rect 485 276 486 277
rect 486 276 487 277
rect 487 276 488 277
rect 488 276 489 277
rect 489 276 490 277
rect 490 276 491 277
rect 491 276 492 277
rect 492 276 493 277
rect 493 276 494 277
rect 494 276 495 277
rect 495 276 496 277
rect 530 276 531 277
rect 531 276 532 277
rect 532 276 533 277
rect 533 276 534 277
rect 534 276 535 277
rect 535 276 536 277
rect 536 276 537 277
rect 537 276 538 277
rect 538 276 539 277
rect 87 275 88 276
rect 88 275 89 276
rect 89 275 90 276
rect 90 275 91 276
rect 91 275 92 276
rect 92 275 93 276
rect 93 275 94 276
rect 94 275 95 276
rect 95 275 96 276
rect 96 275 97 276
rect 97 275 98 276
rect 98 275 99 276
rect 126 275 127 276
rect 127 275 128 276
rect 128 275 129 276
rect 129 275 130 276
rect 130 275 131 276
rect 131 275 132 276
rect 132 275 133 276
rect 133 275 134 276
rect 134 275 135 276
rect 135 275 136 276
rect 141 275 142 276
rect 142 275 143 276
rect 143 275 144 276
rect 144 275 145 276
rect 145 275 146 276
rect 146 275 147 276
rect 147 275 148 276
rect 148 275 149 276
rect 474 275 475 276
rect 475 275 476 276
rect 476 275 477 276
rect 477 275 478 276
rect 478 275 479 276
rect 479 275 480 276
rect 480 275 481 276
rect 481 275 482 276
rect 482 275 483 276
rect 483 275 484 276
rect 484 275 485 276
rect 485 275 486 276
rect 486 275 487 276
rect 487 275 488 276
rect 488 275 489 276
rect 489 275 490 276
rect 530 275 531 276
rect 531 275 532 276
rect 532 275 533 276
rect 533 275 534 276
rect 534 275 535 276
rect 535 275 536 276
rect 536 275 537 276
rect 537 275 538 276
rect 538 275 539 276
rect 87 274 88 275
rect 88 274 89 275
rect 89 274 90 275
rect 90 274 91 275
rect 91 274 92 275
rect 92 274 93 275
rect 93 274 94 275
rect 94 274 95 275
rect 95 274 96 275
rect 96 274 97 275
rect 97 274 98 275
rect 98 274 99 275
rect 126 274 127 275
rect 127 274 128 275
rect 128 274 129 275
rect 129 274 130 275
rect 130 274 131 275
rect 131 274 132 275
rect 132 274 133 275
rect 133 274 134 275
rect 134 274 135 275
rect 135 274 136 275
rect 136 274 137 275
rect 137 274 138 275
rect 139 274 140 275
rect 140 274 141 275
rect 141 274 142 275
rect 142 274 143 275
rect 143 274 144 275
rect 144 274 145 275
rect 145 274 146 275
rect 146 274 147 275
rect 147 274 148 275
rect 148 274 149 275
rect 474 274 475 275
rect 475 274 476 275
rect 476 274 477 275
rect 477 274 478 275
rect 478 274 479 275
rect 479 274 480 275
rect 480 274 481 275
rect 481 274 482 275
rect 482 274 483 275
rect 483 274 484 275
rect 484 274 485 275
rect 485 274 486 275
rect 486 274 487 275
rect 487 274 488 275
rect 488 274 489 275
rect 489 274 490 275
rect 530 274 531 275
rect 531 274 532 275
rect 532 274 533 275
rect 533 274 534 275
rect 534 274 535 275
rect 535 274 536 275
rect 536 274 537 275
rect 537 274 538 275
rect 538 274 539 275
rect 88 273 89 274
rect 89 273 90 274
rect 90 273 91 274
rect 91 273 92 274
rect 92 273 93 274
rect 93 273 94 274
rect 94 273 95 274
rect 95 273 96 274
rect 96 273 97 274
rect 97 273 98 274
rect 98 273 99 274
rect 128 273 129 274
rect 129 273 130 274
rect 130 273 131 274
rect 131 273 132 274
rect 132 273 133 274
rect 133 273 134 274
rect 134 273 135 274
rect 135 273 136 274
rect 136 273 137 274
rect 137 273 138 274
rect 139 273 140 274
rect 140 273 141 274
rect 141 273 142 274
rect 142 273 143 274
rect 143 273 144 274
rect 144 273 145 274
rect 145 273 146 274
rect 146 273 147 274
rect 147 273 148 274
rect 476 273 477 274
rect 477 273 478 274
rect 478 273 479 274
rect 479 273 480 274
rect 480 273 481 274
rect 481 273 482 274
rect 482 273 483 274
rect 483 273 484 274
rect 484 273 485 274
rect 485 273 486 274
rect 486 273 487 274
rect 532 273 533 274
rect 533 273 534 274
rect 534 273 535 274
rect 535 273 536 274
rect 536 273 537 274
rect 537 273 538 274
rect 538 273 539 274
rect 88 272 89 273
rect 89 272 90 273
rect 90 272 91 273
rect 91 272 92 273
rect 92 272 93 273
rect 93 272 94 273
rect 94 272 95 273
rect 95 272 96 273
rect 96 272 97 273
rect 97 272 98 273
rect 98 272 99 273
rect 126 272 127 273
rect 127 272 128 273
rect 128 272 129 273
rect 129 272 130 273
rect 130 272 131 273
rect 131 272 132 273
rect 132 272 133 273
rect 133 272 134 273
rect 134 272 135 273
rect 135 272 136 273
rect 136 272 137 273
rect 137 272 138 273
rect 138 272 139 273
rect 139 272 140 273
rect 140 272 141 273
rect 141 272 142 273
rect 142 272 143 273
rect 143 272 144 273
rect 144 272 145 273
rect 145 272 146 273
rect 146 272 147 273
rect 147 272 148 273
rect 148 272 149 273
rect 476 272 477 273
rect 477 272 478 273
rect 478 272 479 273
rect 479 272 480 273
rect 480 272 481 273
rect 481 272 482 273
rect 482 272 483 273
rect 483 272 484 273
rect 484 272 485 273
rect 485 272 486 273
rect 486 272 487 273
rect 487 272 488 273
rect 530 272 531 273
rect 531 272 532 273
rect 532 272 533 273
rect 533 272 534 273
rect 534 272 535 273
rect 535 272 536 273
rect 536 272 537 273
rect 537 272 538 273
rect 538 272 539 273
rect 88 271 89 272
rect 89 271 90 272
rect 90 271 91 272
rect 91 271 92 272
rect 92 271 93 272
rect 93 271 94 272
rect 94 271 95 272
rect 95 271 96 272
rect 96 271 97 272
rect 97 271 98 272
rect 98 271 99 272
rect 126 271 127 272
rect 127 271 128 272
rect 128 271 129 272
rect 129 271 130 272
rect 130 271 131 272
rect 131 271 132 272
rect 132 271 133 272
rect 133 271 134 272
rect 134 271 135 272
rect 135 271 136 272
rect 136 271 137 272
rect 137 271 138 272
rect 138 271 139 272
rect 139 271 140 272
rect 140 271 141 272
rect 141 271 142 272
rect 142 271 143 272
rect 143 271 144 272
rect 144 271 145 272
rect 145 271 146 272
rect 146 271 147 272
rect 147 271 148 272
rect 148 271 149 272
rect 476 271 477 272
rect 477 271 478 272
rect 478 271 479 272
rect 479 271 480 272
rect 480 271 481 272
rect 481 271 482 272
rect 482 271 483 272
rect 483 271 484 272
rect 484 271 485 272
rect 485 271 486 272
rect 486 271 487 272
rect 487 271 488 272
rect 530 271 531 272
rect 531 271 532 272
rect 532 271 533 272
rect 533 271 534 272
rect 534 271 535 272
rect 535 271 536 272
rect 536 271 537 272
rect 537 271 538 272
rect 538 271 539 272
rect 88 270 89 271
rect 89 270 90 271
rect 90 270 91 271
rect 91 270 92 271
rect 92 270 93 271
rect 93 270 94 271
rect 94 270 95 271
rect 95 270 96 271
rect 96 270 97 271
rect 97 270 98 271
rect 98 270 99 271
rect 126 270 127 271
rect 127 270 128 271
rect 128 270 129 271
rect 129 270 130 271
rect 130 270 131 271
rect 131 270 132 271
rect 132 270 133 271
rect 133 270 134 271
rect 134 270 135 271
rect 135 270 136 271
rect 136 270 137 271
rect 137 270 138 271
rect 138 270 139 271
rect 139 270 140 271
rect 140 270 141 271
rect 141 270 142 271
rect 142 270 143 271
rect 143 270 144 271
rect 144 270 145 271
rect 145 270 146 271
rect 146 270 147 271
rect 147 270 148 271
rect 148 270 149 271
rect 476 270 477 271
rect 477 270 478 271
rect 478 270 479 271
rect 479 270 480 271
rect 480 270 481 271
rect 481 270 482 271
rect 482 270 483 271
rect 483 270 484 271
rect 484 270 485 271
rect 485 270 486 271
rect 486 270 487 271
rect 487 270 488 271
rect 530 270 531 271
rect 531 270 532 271
rect 532 270 533 271
rect 533 270 534 271
rect 534 270 535 271
rect 535 270 536 271
rect 536 270 537 271
rect 537 270 538 271
rect 538 270 539 271
rect 90 269 91 270
rect 91 269 92 270
rect 92 269 93 270
rect 93 269 94 270
rect 94 269 95 270
rect 95 269 96 270
rect 96 269 97 270
rect 97 269 98 270
rect 98 269 99 270
rect 126 269 127 270
rect 127 269 128 270
rect 128 269 129 270
rect 129 269 130 270
rect 130 269 131 270
rect 131 269 132 270
rect 132 269 133 270
rect 133 269 134 270
rect 134 269 135 270
rect 135 269 136 270
rect 136 269 137 270
rect 137 269 138 270
rect 138 269 139 270
rect 139 269 140 270
rect 140 269 141 270
rect 141 269 142 270
rect 142 269 143 270
rect 143 269 144 270
rect 144 269 145 270
rect 145 269 146 270
rect 146 269 147 270
rect 147 269 148 270
rect 148 269 149 270
rect 476 269 477 270
rect 477 269 478 270
rect 478 269 479 270
rect 479 269 480 270
rect 480 269 481 270
rect 481 269 482 270
rect 482 269 483 270
rect 483 269 484 270
rect 484 269 485 270
rect 485 269 486 270
rect 486 269 487 270
rect 487 269 488 270
rect 530 269 531 270
rect 531 269 532 270
rect 532 269 533 270
rect 533 269 534 270
rect 534 269 535 270
rect 535 269 536 270
rect 536 269 537 270
rect 537 269 538 270
rect 538 269 539 270
rect 90 268 91 269
rect 91 268 92 269
rect 92 268 93 269
rect 93 268 94 269
rect 94 268 95 269
rect 95 268 96 269
rect 96 268 97 269
rect 97 268 98 269
rect 98 268 99 269
rect 126 268 127 269
rect 127 268 128 269
rect 128 268 129 269
rect 129 268 130 269
rect 130 268 131 269
rect 131 268 132 269
rect 132 268 133 269
rect 133 268 134 269
rect 134 268 135 269
rect 135 268 136 269
rect 136 268 137 269
rect 137 268 138 269
rect 138 268 139 269
rect 139 268 140 269
rect 140 268 141 269
rect 141 268 142 269
rect 142 268 143 269
rect 143 268 144 269
rect 144 268 145 269
rect 145 268 146 269
rect 146 268 147 269
rect 147 268 148 269
rect 148 268 149 269
rect 149 268 150 269
rect 150 268 151 269
rect 476 268 477 269
rect 477 268 478 269
rect 478 268 479 269
rect 479 268 480 269
rect 480 268 481 269
rect 481 268 482 269
rect 482 268 483 269
rect 483 268 484 269
rect 484 268 485 269
rect 485 268 486 269
rect 486 268 487 269
rect 487 268 488 269
rect 530 268 531 269
rect 531 268 532 269
rect 532 268 533 269
rect 533 268 534 269
rect 534 268 535 269
rect 535 268 536 269
rect 536 268 537 269
rect 537 268 538 269
rect 538 268 539 269
rect 92 267 93 268
rect 93 267 94 268
rect 94 267 95 268
rect 95 267 96 268
rect 96 267 97 268
rect 97 267 98 268
rect 98 267 99 268
rect 126 267 127 268
rect 127 267 128 268
rect 128 267 129 268
rect 129 267 130 268
rect 130 267 131 268
rect 131 267 132 268
rect 132 267 133 268
rect 133 267 134 268
rect 134 267 135 268
rect 135 267 136 268
rect 136 267 137 268
rect 137 267 138 268
rect 138 267 139 268
rect 139 267 140 268
rect 140 267 141 268
rect 141 267 142 268
rect 142 267 143 268
rect 143 267 144 268
rect 144 267 145 268
rect 145 267 146 268
rect 146 267 147 268
rect 147 267 148 268
rect 148 267 149 268
rect 149 267 150 268
rect 150 267 151 268
rect 476 267 477 268
rect 477 267 478 268
rect 478 267 479 268
rect 479 267 480 268
rect 480 267 481 268
rect 481 267 482 268
rect 482 267 483 268
rect 483 267 484 268
rect 484 267 485 268
rect 485 267 486 268
rect 486 267 487 268
rect 487 267 488 268
rect 530 267 531 268
rect 531 267 532 268
rect 532 267 533 268
rect 533 267 534 268
rect 534 267 535 268
rect 535 267 536 268
rect 536 267 537 268
rect 537 267 538 268
rect 538 267 539 268
rect 92 266 93 267
rect 93 266 94 267
rect 94 266 95 267
rect 95 266 96 267
rect 96 266 97 267
rect 97 266 98 267
rect 98 266 99 267
rect 126 266 127 267
rect 127 266 128 267
rect 128 266 129 267
rect 129 266 130 267
rect 130 266 131 267
rect 131 266 132 267
rect 132 266 133 267
rect 133 266 134 267
rect 134 266 135 267
rect 135 266 136 267
rect 136 266 137 267
rect 137 266 138 267
rect 138 266 139 267
rect 139 266 140 267
rect 140 266 141 267
rect 141 266 142 267
rect 142 266 143 267
rect 143 266 144 267
rect 144 266 145 267
rect 145 266 146 267
rect 146 266 147 267
rect 147 266 148 267
rect 148 266 149 267
rect 149 266 150 267
rect 150 266 151 267
rect 151 266 152 267
rect 152 266 153 267
rect 476 266 477 267
rect 477 266 478 267
rect 478 266 479 267
rect 479 266 480 267
rect 480 266 481 267
rect 481 266 482 267
rect 482 266 483 267
rect 483 266 484 267
rect 484 266 485 267
rect 485 266 486 267
rect 486 266 487 267
rect 487 266 488 267
rect 530 266 531 267
rect 531 266 532 267
rect 532 266 533 267
rect 533 266 534 267
rect 534 266 535 267
rect 535 266 536 267
rect 536 266 537 267
rect 537 266 538 267
rect 538 266 539 267
rect 92 265 93 266
rect 93 265 94 266
rect 94 265 95 266
rect 95 265 96 266
rect 96 265 97 266
rect 126 265 127 266
rect 127 265 128 266
rect 128 265 129 266
rect 129 265 130 266
rect 130 265 131 266
rect 131 265 132 266
rect 132 265 133 266
rect 133 265 134 266
rect 134 265 135 266
rect 135 265 136 266
rect 136 265 137 266
rect 137 265 138 266
rect 139 265 140 266
rect 140 265 141 266
rect 141 265 142 266
rect 142 265 143 266
rect 143 265 144 266
rect 144 265 145 266
rect 145 265 146 266
rect 146 265 147 266
rect 147 265 148 266
rect 148 265 149 266
rect 149 265 150 266
rect 150 265 151 266
rect 151 265 152 266
rect 152 265 153 266
rect 476 265 477 266
rect 477 265 478 266
rect 478 265 479 266
rect 479 265 480 266
rect 480 265 481 266
rect 481 265 482 266
rect 482 265 483 266
rect 483 265 484 266
rect 484 265 485 266
rect 485 265 486 266
rect 486 265 487 266
rect 487 265 488 266
rect 532 265 533 266
rect 533 265 534 266
rect 534 265 535 266
rect 535 265 536 266
rect 536 265 537 266
rect 537 265 538 266
rect 538 265 539 266
rect 92 264 93 265
rect 93 264 94 265
rect 94 264 95 265
rect 95 264 96 265
rect 96 264 97 265
rect 126 264 127 265
rect 127 264 128 265
rect 128 264 129 265
rect 129 264 130 265
rect 130 264 131 265
rect 131 264 132 265
rect 132 264 133 265
rect 133 264 134 265
rect 134 264 135 265
rect 135 264 136 265
rect 136 264 137 265
rect 137 264 138 265
rect 139 264 140 265
rect 140 264 141 265
rect 141 264 142 265
rect 142 264 143 265
rect 143 264 144 265
rect 144 264 145 265
rect 145 264 146 265
rect 146 264 147 265
rect 147 264 148 265
rect 148 264 149 265
rect 149 264 150 265
rect 150 264 151 265
rect 151 264 152 265
rect 152 264 153 265
rect 153 264 154 265
rect 154 264 155 265
rect 476 264 477 265
rect 477 264 478 265
rect 478 264 479 265
rect 479 264 480 265
rect 480 264 481 265
rect 481 264 482 265
rect 482 264 483 265
rect 483 264 484 265
rect 484 264 485 265
rect 485 264 486 265
rect 486 264 487 265
rect 487 264 488 265
rect 530 264 531 265
rect 531 264 532 265
rect 532 264 533 265
rect 533 264 534 265
rect 534 264 535 265
rect 535 264 536 265
rect 536 264 537 265
rect 537 264 538 265
rect 538 264 539 265
rect 94 263 95 264
rect 95 263 96 264
rect 96 263 97 264
rect 126 263 127 264
rect 127 263 128 264
rect 128 263 129 264
rect 129 263 130 264
rect 130 263 131 264
rect 131 263 132 264
rect 132 263 133 264
rect 133 263 134 264
rect 134 263 135 264
rect 135 263 136 264
rect 141 263 142 264
rect 142 263 143 264
rect 143 263 144 264
rect 144 263 145 264
rect 145 263 146 264
rect 146 263 147 264
rect 147 263 148 264
rect 148 263 149 264
rect 149 263 150 264
rect 150 263 151 264
rect 151 263 152 264
rect 152 263 153 264
rect 153 263 154 264
rect 154 263 155 264
rect 476 263 477 264
rect 477 263 478 264
rect 478 263 479 264
rect 479 263 480 264
rect 480 263 481 264
rect 481 263 482 264
rect 482 263 483 264
rect 483 263 484 264
rect 484 263 485 264
rect 485 263 486 264
rect 486 263 487 264
rect 530 263 531 264
rect 531 263 532 264
rect 532 263 533 264
rect 533 263 534 264
rect 534 263 535 264
rect 535 263 536 264
rect 536 263 537 264
rect 537 263 538 264
rect 538 263 539 264
rect 94 262 95 263
rect 95 262 96 263
rect 96 262 97 263
rect 126 262 127 263
rect 127 262 128 263
rect 128 262 129 263
rect 129 262 130 263
rect 130 262 131 263
rect 131 262 132 263
rect 132 262 133 263
rect 133 262 134 263
rect 134 262 135 263
rect 135 262 136 263
rect 136 262 137 263
rect 137 262 138 263
rect 141 262 142 263
rect 142 262 143 263
rect 143 262 144 263
rect 144 262 145 263
rect 145 262 146 263
rect 146 262 147 263
rect 147 262 148 263
rect 148 262 149 263
rect 149 262 150 263
rect 150 262 151 263
rect 151 262 152 263
rect 152 262 153 263
rect 153 262 154 263
rect 154 262 155 263
rect 155 262 156 263
rect 156 262 157 263
rect 476 262 477 263
rect 477 262 478 263
rect 478 262 479 263
rect 479 262 480 263
rect 480 262 481 263
rect 481 262 482 263
rect 482 262 483 263
rect 483 262 484 263
rect 484 262 485 263
rect 485 262 486 263
rect 486 262 487 263
rect 487 262 488 263
rect 530 262 531 263
rect 531 262 532 263
rect 532 262 533 263
rect 533 262 534 263
rect 534 262 535 263
rect 535 262 536 263
rect 536 262 537 263
rect 537 262 538 263
rect 538 262 539 263
rect 94 261 95 262
rect 95 261 96 262
rect 96 261 97 262
rect 126 261 127 262
rect 127 261 128 262
rect 128 261 129 262
rect 129 261 130 262
rect 130 261 131 262
rect 131 261 132 262
rect 132 261 133 262
rect 133 261 134 262
rect 134 261 135 262
rect 135 261 136 262
rect 136 261 137 262
rect 137 261 138 262
rect 143 261 144 262
rect 144 261 145 262
rect 145 261 146 262
rect 146 261 147 262
rect 147 261 148 262
rect 148 261 149 262
rect 149 261 150 262
rect 150 261 151 262
rect 151 261 152 262
rect 152 261 153 262
rect 153 261 154 262
rect 154 261 155 262
rect 155 261 156 262
rect 156 261 157 262
rect 476 261 477 262
rect 477 261 478 262
rect 478 261 479 262
rect 479 261 480 262
rect 480 261 481 262
rect 481 261 482 262
rect 482 261 483 262
rect 483 261 484 262
rect 484 261 485 262
rect 485 261 486 262
rect 486 261 487 262
rect 487 261 488 262
rect 530 261 531 262
rect 531 261 532 262
rect 532 261 533 262
rect 533 261 534 262
rect 534 261 535 262
rect 535 261 536 262
rect 536 261 537 262
rect 537 261 538 262
rect 538 261 539 262
rect 94 260 95 261
rect 95 260 96 261
rect 96 260 97 261
rect 126 260 127 261
rect 127 260 128 261
rect 128 260 129 261
rect 129 260 130 261
rect 130 260 131 261
rect 131 260 132 261
rect 132 260 133 261
rect 133 260 134 261
rect 134 260 135 261
rect 135 260 136 261
rect 136 260 137 261
rect 137 260 138 261
rect 143 260 144 261
rect 144 260 145 261
rect 145 260 146 261
rect 146 260 147 261
rect 147 260 148 261
rect 148 260 149 261
rect 149 260 150 261
rect 150 260 151 261
rect 151 260 152 261
rect 152 260 153 261
rect 153 260 154 261
rect 154 260 155 261
rect 155 260 156 261
rect 156 260 157 261
rect 157 260 158 261
rect 158 260 159 261
rect 191 260 192 261
rect 192 260 193 261
rect 193 260 194 261
rect 194 260 195 261
rect 195 260 196 261
rect 476 260 477 261
rect 477 260 478 261
rect 478 260 479 261
rect 479 260 480 261
rect 480 260 481 261
rect 481 260 482 261
rect 482 260 483 261
rect 483 260 484 261
rect 484 260 485 261
rect 485 260 486 261
rect 486 260 487 261
rect 487 260 488 261
rect 530 260 531 261
rect 531 260 532 261
rect 532 260 533 261
rect 533 260 534 261
rect 534 260 535 261
rect 535 260 536 261
rect 536 260 537 261
rect 537 260 538 261
rect 538 260 539 261
rect 94 259 95 260
rect 95 259 96 260
rect 96 259 97 260
rect 126 259 127 260
rect 127 259 128 260
rect 128 259 129 260
rect 129 259 130 260
rect 130 259 131 260
rect 131 259 132 260
rect 132 259 133 260
rect 133 259 134 260
rect 134 259 135 260
rect 135 259 136 260
rect 136 259 137 260
rect 137 259 138 260
rect 145 259 146 260
rect 146 259 147 260
rect 147 259 148 260
rect 148 259 149 260
rect 149 259 150 260
rect 150 259 151 260
rect 151 259 152 260
rect 152 259 153 260
rect 153 259 154 260
rect 154 259 155 260
rect 155 259 156 260
rect 156 259 157 260
rect 157 259 158 260
rect 158 259 159 260
rect 191 259 192 260
rect 192 259 193 260
rect 193 259 194 260
rect 194 259 195 260
rect 195 259 196 260
rect 476 259 477 260
rect 477 259 478 260
rect 478 259 479 260
rect 479 259 480 260
rect 480 259 481 260
rect 481 259 482 260
rect 482 259 483 260
rect 483 259 484 260
rect 484 259 485 260
rect 485 259 486 260
rect 486 259 487 260
rect 487 259 488 260
rect 530 259 531 260
rect 531 259 532 260
rect 532 259 533 260
rect 533 259 534 260
rect 534 259 535 260
rect 535 259 536 260
rect 536 259 537 260
rect 537 259 538 260
rect 538 259 539 260
rect 94 258 95 259
rect 95 258 96 259
rect 96 258 97 259
rect 126 258 127 259
rect 127 258 128 259
rect 128 258 129 259
rect 129 258 130 259
rect 130 258 131 259
rect 131 258 132 259
rect 132 258 133 259
rect 133 258 134 259
rect 134 258 135 259
rect 135 258 136 259
rect 136 258 137 259
rect 137 258 138 259
rect 145 258 146 259
rect 146 258 147 259
rect 147 258 148 259
rect 148 258 149 259
rect 149 258 150 259
rect 150 258 151 259
rect 151 258 152 259
rect 152 258 153 259
rect 153 258 154 259
rect 154 258 155 259
rect 155 258 156 259
rect 156 258 157 259
rect 157 258 158 259
rect 158 258 159 259
rect 159 258 160 259
rect 160 258 161 259
rect 191 258 192 259
rect 192 258 193 259
rect 193 258 194 259
rect 194 258 195 259
rect 195 258 196 259
rect 196 258 197 259
rect 197 258 198 259
rect 476 258 477 259
rect 477 258 478 259
rect 478 258 479 259
rect 479 258 480 259
rect 480 258 481 259
rect 481 258 482 259
rect 482 258 483 259
rect 483 258 484 259
rect 484 258 485 259
rect 485 258 486 259
rect 486 258 487 259
rect 487 258 488 259
rect 530 258 531 259
rect 531 258 532 259
rect 532 258 533 259
rect 533 258 534 259
rect 534 258 535 259
rect 535 258 536 259
rect 536 258 537 259
rect 537 258 538 259
rect 538 258 539 259
rect 126 257 127 258
rect 127 257 128 258
rect 128 257 129 258
rect 129 257 130 258
rect 130 257 131 258
rect 131 257 132 258
rect 132 257 133 258
rect 133 257 134 258
rect 134 257 135 258
rect 135 257 136 258
rect 136 257 137 258
rect 137 257 138 258
rect 147 257 148 258
rect 148 257 149 258
rect 149 257 150 258
rect 150 257 151 258
rect 151 257 152 258
rect 152 257 153 258
rect 153 257 154 258
rect 154 257 155 258
rect 155 257 156 258
rect 156 257 157 258
rect 157 257 158 258
rect 158 257 159 258
rect 159 257 160 258
rect 160 257 161 258
rect 191 257 192 258
rect 192 257 193 258
rect 193 257 194 258
rect 194 257 195 258
rect 195 257 196 258
rect 196 257 197 258
rect 197 257 198 258
rect 476 257 477 258
rect 477 257 478 258
rect 478 257 479 258
rect 479 257 480 258
rect 480 257 481 258
rect 481 257 482 258
rect 482 257 483 258
rect 483 257 484 258
rect 484 257 485 258
rect 485 257 486 258
rect 486 257 487 258
rect 532 257 533 258
rect 533 257 534 258
rect 534 257 535 258
rect 535 257 536 258
rect 536 257 537 258
rect 537 257 538 258
rect 538 257 539 258
rect 126 256 127 257
rect 127 256 128 257
rect 128 256 129 257
rect 129 256 130 257
rect 130 256 131 257
rect 131 256 132 257
rect 132 256 133 257
rect 133 256 134 257
rect 134 256 135 257
rect 135 256 136 257
rect 136 256 137 257
rect 137 256 138 257
rect 147 256 148 257
rect 148 256 149 257
rect 149 256 150 257
rect 150 256 151 257
rect 151 256 152 257
rect 152 256 153 257
rect 153 256 154 257
rect 154 256 155 257
rect 155 256 156 257
rect 156 256 157 257
rect 157 256 158 257
rect 158 256 159 257
rect 159 256 160 257
rect 160 256 161 257
rect 190 256 191 257
rect 191 256 192 257
rect 192 256 193 257
rect 193 256 194 257
rect 194 256 195 257
rect 195 256 196 257
rect 196 256 197 257
rect 197 256 198 257
rect 476 256 477 257
rect 477 256 478 257
rect 478 256 479 257
rect 479 256 480 257
rect 480 256 481 257
rect 481 256 482 257
rect 482 256 483 257
rect 483 256 484 257
rect 484 256 485 257
rect 485 256 486 257
rect 486 256 487 257
rect 487 256 488 257
rect 530 256 531 257
rect 531 256 532 257
rect 532 256 533 257
rect 533 256 534 257
rect 534 256 535 257
rect 535 256 536 257
rect 536 256 537 257
rect 537 256 538 257
rect 538 256 539 257
rect 126 255 127 256
rect 127 255 128 256
rect 128 255 129 256
rect 129 255 130 256
rect 130 255 131 256
rect 131 255 132 256
rect 132 255 133 256
rect 133 255 134 256
rect 134 255 135 256
rect 135 255 136 256
rect 148 255 149 256
rect 149 255 150 256
rect 150 255 151 256
rect 151 255 152 256
rect 152 255 153 256
rect 153 255 154 256
rect 154 255 155 256
rect 155 255 156 256
rect 156 255 157 256
rect 157 255 158 256
rect 158 255 159 256
rect 159 255 160 256
rect 160 255 161 256
rect 190 255 191 256
rect 191 255 192 256
rect 192 255 193 256
rect 193 255 194 256
rect 194 255 195 256
rect 195 255 196 256
rect 196 255 197 256
rect 197 255 198 256
rect 476 255 477 256
rect 477 255 478 256
rect 478 255 479 256
rect 479 255 480 256
rect 480 255 481 256
rect 481 255 482 256
rect 482 255 483 256
rect 483 255 484 256
rect 484 255 485 256
rect 485 255 486 256
rect 486 255 487 256
rect 487 255 488 256
rect 530 255 531 256
rect 531 255 532 256
rect 532 255 533 256
rect 533 255 534 256
rect 534 255 535 256
rect 535 255 536 256
rect 536 255 537 256
rect 537 255 538 256
rect 538 255 539 256
rect 94 254 95 255
rect 95 254 96 255
rect 96 254 97 255
rect 126 254 127 255
rect 127 254 128 255
rect 128 254 129 255
rect 129 254 130 255
rect 130 254 131 255
rect 131 254 132 255
rect 132 254 133 255
rect 133 254 134 255
rect 134 254 135 255
rect 135 254 136 255
rect 136 254 137 255
rect 137 254 138 255
rect 148 254 149 255
rect 149 254 150 255
rect 150 254 151 255
rect 151 254 152 255
rect 152 254 153 255
rect 153 254 154 255
rect 154 254 155 255
rect 155 254 156 255
rect 156 254 157 255
rect 157 254 158 255
rect 158 254 159 255
rect 159 254 160 255
rect 160 254 161 255
rect 161 254 162 255
rect 162 254 163 255
rect 163 254 164 255
rect 190 254 191 255
rect 191 254 192 255
rect 192 254 193 255
rect 193 254 194 255
rect 194 254 195 255
rect 195 254 196 255
rect 196 254 197 255
rect 197 254 198 255
rect 476 254 477 255
rect 477 254 478 255
rect 478 254 479 255
rect 479 254 480 255
rect 480 254 481 255
rect 481 254 482 255
rect 482 254 483 255
rect 483 254 484 255
rect 484 254 485 255
rect 485 254 486 255
rect 486 254 487 255
rect 487 254 488 255
rect 530 254 531 255
rect 531 254 532 255
rect 532 254 533 255
rect 533 254 534 255
rect 534 254 535 255
rect 535 254 536 255
rect 536 254 537 255
rect 537 254 538 255
rect 538 254 539 255
rect 94 253 95 254
rect 95 253 96 254
rect 96 253 97 254
rect 128 253 129 254
rect 129 253 130 254
rect 130 253 131 254
rect 131 253 132 254
rect 132 253 133 254
rect 133 253 134 254
rect 134 253 135 254
rect 135 253 136 254
rect 136 253 137 254
rect 137 253 138 254
rect 150 253 151 254
rect 151 253 152 254
rect 152 253 153 254
rect 153 253 154 254
rect 154 253 155 254
rect 155 253 156 254
rect 156 253 157 254
rect 157 253 158 254
rect 158 253 159 254
rect 159 253 160 254
rect 160 253 161 254
rect 161 253 162 254
rect 162 253 163 254
rect 163 253 164 254
rect 190 253 191 254
rect 191 253 192 254
rect 192 253 193 254
rect 193 253 194 254
rect 194 253 195 254
rect 195 253 196 254
rect 196 253 197 254
rect 197 253 198 254
rect 476 253 477 254
rect 477 253 478 254
rect 478 253 479 254
rect 479 253 480 254
rect 480 253 481 254
rect 481 253 482 254
rect 482 253 483 254
rect 483 253 484 254
rect 484 253 485 254
rect 485 253 486 254
rect 486 253 487 254
rect 487 253 488 254
rect 530 253 531 254
rect 531 253 532 254
rect 532 253 533 254
rect 533 253 534 254
rect 534 253 535 254
rect 535 253 536 254
rect 536 253 537 254
rect 537 253 538 254
rect 538 253 539 254
rect 94 252 95 253
rect 95 252 96 253
rect 96 252 97 253
rect 126 252 127 253
rect 127 252 128 253
rect 128 252 129 253
rect 129 252 130 253
rect 130 252 131 253
rect 131 252 132 253
rect 132 252 133 253
rect 133 252 134 253
rect 134 252 135 253
rect 135 252 136 253
rect 136 252 137 253
rect 137 252 138 253
rect 150 252 151 253
rect 151 252 152 253
rect 152 252 153 253
rect 153 252 154 253
rect 154 252 155 253
rect 155 252 156 253
rect 156 252 157 253
rect 157 252 158 253
rect 158 252 159 253
rect 159 252 160 253
rect 160 252 161 253
rect 161 252 162 253
rect 162 252 163 253
rect 163 252 164 253
rect 164 252 165 253
rect 165 252 166 253
rect 188 252 189 253
rect 189 252 190 253
rect 190 252 191 253
rect 191 252 192 253
rect 192 252 193 253
rect 193 252 194 253
rect 194 252 195 253
rect 195 252 196 253
rect 196 252 197 253
rect 197 252 198 253
rect 198 252 199 253
rect 199 252 200 253
rect 476 252 477 253
rect 477 252 478 253
rect 478 252 479 253
rect 479 252 480 253
rect 480 252 481 253
rect 481 252 482 253
rect 482 252 483 253
rect 483 252 484 253
rect 484 252 485 253
rect 485 252 486 253
rect 486 252 487 253
rect 487 252 488 253
rect 530 252 531 253
rect 531 252 532 253
rect 532 252 533 253
rect 533 252 534 253
rect 534 252 535 253
rect 535 252 536 253
rect 536 252 537 253
rect 537 252 538 253
rect 538 252 539 253
rect 94 251 95 252
rect 95 251 96 252
rect 96 251 97 252
rect 126 251 127 252
rect 127 251 128 252
rect 128 251 129 252
rect 129 251 130 252
rect 130 251 131 252
rect 131 251 132 252
rect 132 251 133 252
rect 133 251 134 252
rect 134 251 135 252
rect 135 251 136 252
rect 136 251 137 252
rect 137 251 138 252
rect 152 251 153 252
rect 153 251 154 252
rect 154 251 155 252
rect 155 251 156 252
rect 156 251 157 252
rect 157 251 158 252
rect 158 251 159 252
rect 159 251 160 252
rect 160 251 161 252
rect 161 251 162 252
rect 162 251 163 252
rect 163 251 164 252
rect 164 251 165 252
rect 165 251 166 252
rect 188 251 189 252
rect 189 251 190 252
rect 190 251 191 252
rect 191 251 192 252
rect 192 251 193 252
rect 193 251 194 252
rect 194 251 195 252
rect 195 251 196 252
rect 196 251 197 252
rect 197 251 198 252
rect 198 251 199 252
rect 199 251 200 252
rect 476 251 477 252
rect 477 251 478 252
rect 478 251 479 252
rect 479 251 480 252
rect 480 251 481 252
rect 481 251 482 252
rect 482 251 483 252
rect 483 251 484 252
rect 484 251 485 252
rect 485 251 486 252
rect 486 251 487 252
rect 487 251 488 252
rect 530 251 531 252
rect 531 251 532 252
rect 532 251 533 252
rect 533 251 534 252
rect 534 251 535 252
rect 535 251 536 252
rect 536 251 537 252
rect 537 251 538 252
rect 538 251 539 252
rect 94 250 95 251
rect 95 250 96 251
rect 96 250 97 251
rect 126 250 127 251
rect 127 250 128 251
rect 128 250 129 251
rect 129 250 130 251
rect 130 250 131 251
rect 131 250 132 251
rect 132 250 133 251
rect 133 250 134 251
rect 134 250 135 251
rect 135 250 136 251
rect 136 250 137 251
rect 137 250 138 251
rect 152 250 153 251
rect 153 250 154 251
rect 154 250 155 251
rect 155 250 156 251
rect 156 250 157 251
rect 157 250 158 251
rect 158 250 159 251
rect 159 250 160 251
rect 160 250 161 251
rect 161 250 162 251
rect 162 250 163 251
rect 163 250 164 251
rect 164 250 165 251
rect 165 250 166 251
rect 188 250 189 251
rect 189 250 190 251
rect 190 250 191 251
rect 191 250 192 251
rect 192 250 193 251
rect 193 250 194 251
rect 194 250 195 251
rect 195 250 196 251
rect 196 250 197 251
rect 197 250 198 251
rect 198 250 199 251
rect 199 250 200 251
rect 476 250 477 251
rect 477 250 478 251
rect 478 250 479 251
rect 479 250 480 251
rect 480 250 481 251
rect 481 250 482 251
rect 482 250 483 251
rect 483 250 484 251
rect 484 250 485 251
rect 485 250 486 251
rect 486 250 487 251
rect 487 250 488 251
rect 530 250 531 251
rect 531 250 532 251
rect 532 250 533 251
rect 533 250 534 251
rect 534 250 535 251
rect 535 250 536 251
rect 536 250 537 251
rect 537 250 538 251
rect 538 250 539 251
rect 94 249 95 250
rect 95 249 96 250
rect 96 249 97 250
rect 126 249 127 250
rect 127 249 128 250
rect 128 249 129 250
rect 129 249 130 250
rect 130 249 131 250
rect 131 249 132 250
rect 132 249 133 250
rect 133 249 134 250
rect 134 249 135 250
rect 135 249 136 250
rect 152 249 153 250
rect 153 249 154 250
rect 154 249 155 250
rect 155 249 156 250
rect 156 249 157 250
rect 157 249 158 250
rect 158 249 159 250
rect 159 249 160 250
rect 160 249 161 250
rect 161 249 162 250
rect 162 249 163 250
rect 163 249 164 250
rect 164 249 165 250
rect 165 249 166 250
rect 188 249 189 250
rect 189 249 190 250
rect 190 249 191 250
rect 191 249 192 250
rect 192 249 193 250
rect 193 249 194 250
rect 194 249 195 250
rect 195 249 196 250
rect 196 249 197 250
rect 197 249 198 250
rect 198 249 199 250
rect 199 249 200 250
rect 476 249 477 250
rect 477 249 478 250
rect 478 249 479 250
rect 479 249 480 250
rect 480 249 481 250
rect 481 249 482 250
rect 482 249 483 250
rect 483 249 484 250
rect 484 249 485 250
rect 485 249 486 250
rect 486 249 487 250
rect 487 249 488 250
rect 530 249 531 250
rect 531 249 532 250
rect 532 249 533 250
rect 533 249 534 250
rect 534 249 535 250
rect 535 249 536 250
rect 536 249 537 250
rect 537 249 538 250
rect 538 249 539 250
rect 94 248 95 249
rect 95 248 96 249
rect 96 248 97 249
rect 126 248 127 249
rect 127 248 128 249
rect 128 248 129 249
rect 129 248 130 249
rect 130 248 131 249
rect 131 248 132 249
rect 132 248 133 249
rect 133 248 134 249
rect 134 248 135 249
rect 135 248 136 249
rect 152 248 153 249
rect 153 248 154 249
rect 154 248 155 249
rect 155 248 156 249
rect 156 248 157 249
rect 157 248 158 249
rect 158 248 159 249
rect 159 248 160 249
rect 160 248 161 249
rect 161 248 162 249
rect 162 248 163 249
rect 163 248 164 249
rect 164 248 165 249
rect 165 248 166 249
rect 166 248 167 249
rect 167 248 168 249
rect 188 248 189 249
rect 189 248 190 249
rect 190 248 191 249
rect 191 248 192 249
rect 192 248 193 249
rect 193 248 194 249
rect 194 248 195 249
rect 195 248 196 249
rect 196 248 197 249
rect 197 248 198 249
rect 198 248 199 249
rect 199 248 200 249
rect 200 248 201 249
rect 201 248 202 249
rect 476 248 477 249
rect 477 248 478 249
rect 478 248 479 249
rect 479 248 480 249
rect 480 248 481 249
rect 481 248 482 249
rect 482 248 483 249
rect 483 248 484 249
rect 484 248 485 249
rect 485 248 486 249
rect 486 248 487 249
rect 487 248 488 249
rect 530 248 531 249
rect 531 248 532 249
rect 532 248 533 249
rect 533 248 534 249
rect 534 248 535 249
rect 535 248 536 249
rect 536 248 537 249
rect 537 248 538 249
rect 538 248 539 249
rect 126 247 127 248
rect 127 247 128 248
rect 128 247 129 248
rect 129 247 130 248
rect 130 247 131 248
rect 131 247 132 248
rect 132 247 133 248
rect 133 247 134 248
rect 134 247 135 248
rect 135 247 136 248
rect 154 247 155 248
rect 155 247 156 248
rect 156 247 157 248
rect 157 247 158 248
rect 158 247 159 248
rect 159 247 160 248
rect 160 247 161 248
rect 161 247 162 248
rect 162 247 163 248
rect 163 247 164 248
rect 164 247 165 248
rect 165 247 166 248
rect 166 247 167 248
rect 167 247 168 248
rect 188 247 189 248
rect 189 247 190 248
rect 190 247 191 248
rect 191 247 192 248
rect 192 247 193 248
rect 193 247 194 248
rect 194 247 195 248
rect 195 247 196 248
rect 196 247 197 248
rect 197 247 198 248
rect 198 247 199 248
rect 199 247 200 248
rect 200 247 201 248
rect 201 247 202 248
rect 476 247 477 248
rect 477 247 478 248
rect 478 247 479 248
rect 479 247 480 248
rect 480 247 481 248
rect 481 247 482 248
rect 482 247 483 248
rect 483 247 484 248
rect 484 247 485 248
rect 485 247 486 248
rect 486 247 487 248
rect 530 247 531 248
rect 531 247 532 248
rect 532 247 533 248
rect 533 247 534 248
rect 534 247 535 248
rect 535 247 536 248
rect 536 247 537 248
rect 537 247 538 248
rect 538 247 539 248
rect 94 246 95 247
rect 95 246 96 247
rect 96 246 97 247
rect 126 246 127 247
rect 127 246 128 247
rect 128 246 129 247
rect 129 246 130 247
rect 130 246 131 247
rect 131 246 132 247
rect 132 246 133 247
rect 133 246 134 247
rect 134 246 135 247
rect 135 246 136 247
rect 136 246 137 247
rect 137 246 138 247
rect 154 246 155 247
rect 155 246 156 247
rect 156 246 157 247
rect 157 246 158 247
rect 158 246 159 247
rect 159 246 160 247
rect 160 246 161 247
rect 161 246 162 247
rect 162 246 163 247
rect 163 246 164 247
rect 164 246 165 247
rect 165 246 166 247
rect 166 246 167 247
rect 167 246 168 247
rect 168 246 169 247
rect 169 246 170 247
rect 186 246 187 247
rect 187 246 188 247
rect 188 246 189 247
rect 189 246 190 247
rect 190 246 191 247
rect 191 246 192 247
rect 192 246 193 247
rect 193 246 194 247
rect 194 246 195 247
rect 195 246 196 247
rect 196 246 197 247
rect 197 246 198 247
rect 198 246 199 247
rect 199 246 200 247
rect 200 246 201 247
rect 201 246 202 247
rect 476 246 477 247
rect 477 246 478 247
rect 478 246 479 247
rect 479 246 480 247
rect 480 246 481 247
rect 481 246 482 247
rect 482 246 483 247
rect 483 246 484 247
rect 484 246 485 247
rect 485 246 486 247
rect 486 246 487 247
rect 487 246 488 247
rect 530 246 531 247
rect 531 246 532 247
rect 532 246 533 247
rect 533 246 534 247
rect 534 246 535 247
rect 535 246 536 247
rect 536 246 537 247
rect 537 246 538 247
rect 538 246 539 247
rect 94 245 95 246
rect 95 245 96 246
rect 96 245 97 246
rect 126 245 127 246
rect 127 245 128 246
rect 128 245 129 246
rect 129 245 130 246
rect 130 245 131 246
rect 131 245 132 246
rect 132 245 133 246
rect 133 245 134 246
rect 134 245 135 246
rect 135 245 136 246
rect 136 245 137 246
rect 137 245 138 246
rect 156 245 157 246
rect 157 245 158 246
rect 158 245 159 246
rect 159 245 160 246
rect 160 245 161 246
rect 161 245 162 246
rect 162 245 163 246
rect 163 245 164 246
rect 164 245 165 246
rect 165 245 166 246
rect 166 245 167 246
rect 167 245 168 246
rect 168 245 169 246
rect 169 245 170 246
rect 186 245 187 246
rect 187 245 188 246
rect 188 245 189 246
rect 189 245 190 246
rect 190 245 191 246
rect 191 245 192 246
rect 192 245 193 246
rect 193 245 194 246
rect 194 245 195 246
rect 195 245 196 246
rect 196 245 197 246
rect 197 245 198 246
rect 198 245 199 246
rect 199 245 200 246
rect 200 245 201 246
rect 201 245 202 246
rect 476 245 477 246
rect 477 245 478 246
rect 478 245 479 246
rect 479 245 480 246
rect 480 245 481 246
rect 481 245 482 246
rect 482 245 483 246
rect 483 245 484 246
rect 484 245 485 246
rect 485 245 486 246
rect 486 245 487 246
rect 487 245 488 246
rect 530 245 531 246
rect 531 245 532 246
rect 532 245 533 246
rect 533 245 534 246
rect 534 245 535 246
rect 535 245 536 246
rect 536 245 537 246
rect 94 244 95 245
rect 95 244 96 245
rect 96 244 97 245
rect 126 244 127 245
rect 127 244 128 245
rect 128 244 129 245
rect 129 244 130 245
rect 130 244 131 245
rect 131 244 132 245
rect 132 244 133 245
rect 133 244 134 245
rect 134 244 135 245
rect 135 244 136 245
rect 136 244 137 245
rect 137 244 138 245
rect 156 244 157 245
rect 157 244 158 245
rect 158 244 159 245
rect 159 244 160 245
rect 160 244 161 245
rect 161 244 162 245
rect 162 244 163 245
rect 163 244 164 245
rect 164 244 165 245
rect 165 244 166 245
rect 166 244 167 245
rect 167 244 168 245
rect 168 244 169 245
rect 169 244 170 245
rect 170 244 171 245
rect 171 244 172 245
rect 186 244 187 245
rect 187 244 188 245
rect 188 244 189 245
rect 189 244 190 245
rect 190 244 191 245
rect 191 244 192 245
rect 192 244 193 245
rect 193 244 194 245
rect 194 244 195 245
rect 195 244 196 245
rect 196 244 197 245
rect 197 244 198 245
rect 198 244 199 245
rect 199 244 200 245
rect 200 244 201 245
rect 201 244 202 245
rect 202 244 203 245
rect 203 244 204 245
rect 476 244 477 245
rect 477 244 478 245
rect 478 244 479 245
rect 479 244 480 245
rect 480 244 481 245
rect 481 244 482 245
rect 482 244 483 245
rect 483 244 484 245
rect 484 244 485 245
rect 485 244 486 245
rect 486 244 487 245
rect 487 244 488 245
rect 529 244 530 245
rect 530 244 531 245
rect 531 244 532 245
rect 532 244 533 245
rect 533 244 534 245
rect 534 244 535 245
rect 535 244 536 245
rect 536 244 537 245
rect 126 243 127 244
rect 127 243 128 244
rect 128 243 129 244
rect 129 243 130 244
rect 130 243 131 244
rect 131 243 132 244
rect 132 243 133 244
rect 133 243 134 244
rect 134 243 135 244
rect 135 243 136 244
rect 158 243 159 244
rect 159 243 160 244
rect 160 243 161 244
rect 161 243 162 244
rect 162 243 163 244
rect 163 243 164 244
rect 164 243 165 244
rect 165 243 166 244
rect 166 243 167 244
rect 167 243 168 244
rect 168 243 169 244
rect 169 243 170 244
rect 170 243 171 244
rect 171 243 172 244
rect 186 243 187 244
rect 187 243 188 244
rect 188 243 189 244
rect 189 243 190 244
rect 190 243 191 244
rect 191 243 192 244
rect 192 243 193 244
rect 193 243 194 244
rect 194 243 195 244
rect 195 243 196 244
rect 196 243 197 244
rect 197 243 198 244
rect 198 243 199 244
rect 199 243 200 244
rect 200 243 201 244
rect 201 243 202 244
rect 202 243 203 244
rect 203 243 204 244
rect 476 243 477 244
rect 477 243 478 244
rect 478 243 479 244
rect 479 243 480 244
rect 480 243 481 244
rect 481 243 482 244
rect 482 243 483 244
rect 483 243 484 244
rect 484 243 485 244
rect 485 243 486 244
rect 486 243 487 244
rect 487 243 488 244
rect 529 243 530 244
rect 530 243 531 244
rect 531 243 532 244
rect 532 243 533 244
rect 533 243 534 244
rect 534 243 535 244
rect 535 243 536 244
rect 536 243 537 244
rect 94 242 95 243
rect 95 242 96 243
rect 96 242 97 243
rect 126 242 127 243
rect 127 242 128 243
rect 128 242 129 243
rect 129 242 130 243
rect 130 242 131 243
rect 131 242 132 243
rect 132 242 133 243
rect 133 242 134 243
rect 134 242 135 243
rect 135 242 136 243
rect 136 242 137 243
rect 137 242 138 243
rect 158 242 159 243
rect 159 242 160 243
rect 160 242 161 243
rect 161 242 162 243
rect 162 242 163 243
rect 163 242 164 243
rect 164 242 165 243
rect 165 242 166 243
rect 166 242 167 243
rect 167 242 168 243
rect 168 242 169 243
rect 169 242 170 243
rect 170 242 171 243
rect 171 242 172 243
rect 172 242 173 243
rect 173 242 174 243
rect 184 242 185 243
rect 185 242 186 243
rect 186 242 187 243
rect 187 242 188 243
rect 188 242 189 243
rect 189 242 190 243
rect 190 242 191 243
rect 191 242 192 243
rect 192 242 193 243
rect 193 242 194 243
rect 194 242 195 243
rect 195 242 196 243
rect 196 242 197 243
rect 197 242 198 243
rect 198 242 199 243
rect 199 242 200 243
rect 200 242 201 243
rect 201 242 202 243
rect 202 242 203 243
rect 203 242 204 243
rect 476 242 477 243
rect 477 242 478 243
rect 478 242 479 243
rect 479 242 480 243
rect 480 242 481 243
rect 481 242 482 243
rect 482 242 483 243
rect 483 242 484 243
rect 484 242 485 243
rect 485 242 486 243
rect 486 242 487 243
rect 487 242 488 243
rect 529 242 530 243
rect 530 242 531 243
rect 531 242 532 243
rect 532 242 533 243
rect 533 242 534 243
rect 534 242 535 243
rect 535 242 536 243
rect 536 242 537 243
rect 94 241 95 242
rect 95 241 96 242
rect 96 241 97 242
rect 126 241 127 242
rect 127 241 128 242
rect 128 241 129 242
rect 129 241 130 242
rect 130 241 131 242
rect 131 241 132 242
rect 132 241 133 242
rect 133 241 134 242
rect 134 241 135 242
rect 135 241 136 242
rect 136 241 137 242
rect 137 241 138 242
rect 160 241 161 242
rect 161 241 162 242
rect 162 241 163 242
rect 163 241 164 242
rect 164 241 165 242
rect 165 241 166 242
rect 166 241 167 242
rect 167 241 168 242
rect 168 241 169 242
rect 169 241 170 242
rect 170 241 171 242
rect 171 241 172 242
rect 172 241 173 242
rect 173 241 174 242
rect 184 241 185 242
rect 185 241 186 242
rect 186 241 187 242
rect 187 241 188 242
rect 188 241 189 242
rect 189 241 190 242
rect 190 241 191 242
rect 193 241 194 242
rect 194 241 195 242
rect 195 241 196 242
rect 196 241 197 242
rect 197 241 198 242
rect 198 241 199 242
rect 199 241 200 242
rect 200 241 201 242
rect 201 241 202 242
rect 202 241 203 242
rect 203 241 204 242
rect 476 241 477 242
rect 477 241 478 242
rect 478 241 479 242
rect 479 241 480 242
rect 480 241 481 242
rect 481 241 482 242
rect 482 241 483 242
rect 483 241 484 242
rect 484 241 485 242
rect 485 241 486 242
rect 486 241 487 242
rect 529 241 530 242
rect 530 241 531 242
rect 531 241 532 242
rect 532 241 533 242
rect 533 241 534 242
rect 534 241 535 242
rect 535 241 536 242
rect 536 241 537 242
rect 94 240 95 241
rect 95 240 96 241
rect 96 240 97 241
rect 126 240 127 241
rect 127 240 128 241
rect 128 240 129 241
rect 129 240 130 241
rect 130 240 131 241
rect 131 240 132 241
rect 132 240 133 241
rect 133 240 134 241
rect 134 240 135 241
rect 135 240 136 241
rect 136 240 137 241
rect 137 240 138 241
rect 160 240 161 241
rect 161 240 162 241
rect 162 240 163 241
rect 163 240 164 241
rect 164 240 165 241
rect 165 240 166 241
rect 166 240 167 241
rect 167 240 168 241
rect 168 240 169 241
rect 169 240 170 241
rect 170 240 171 241
rect 171 240 172 241
rect 172 240 173 241
rect 173 240 174 241
rect 174 240 175 241
rect 175 240 176 241
rect 184 240 185 241
rect 185 240 186 241
rect 186 240 187 241
rect 187 240 188 241
rect 188 240 189 241
rect 189 240 190 241
rect 190 240 191 241
rect 193 240 194 241
rect 194 240 195 241
rect 195 240 196 241
rect 196 240 197 241
rect 197 240 198 241
rect 198 240 199 241
rect 199 240 200 241
rect 200 240 201 241
rect 201 240 202 241
rect 202 240 203 241
rect 203 240 204 241
rect 476 240 477 241
rect 477 240 478 241
rect 478 240 479 241
rect 479 240 480 241
rect 480 240 481 241
rect 481 240 482 241
rect 482 240 483 241
rect 483 240 484 241
rect 484 240 485 241
rect 485 240 486 241
rect 486 240 487 241
rect 487 240 488 241
rect 529 240 530 241
rect 530 240 531 241
rect 531 240 532 241
rect 532 240 533 241
rect 533 240 534 241
rect 534 240 535 241
rect 535 240 536 241
rect 536 240 537 241
rect 126 239 127 240
rect 127 239 128 240
rect 128 239 129 240
rect 129 239 130 240
rect 130 239 131 240
rect 131 239 132 240
rect 132 239 133 240
rect 133 239 134 240
rect 134 239 135 240
rect 135 239 136 240
rect 136 239 137 240
rect 137 239 138 240
rect 160 239 161 240
rect 161 239 162 240
rect 162 239 163 240
rect 163 239 164 240
rect 164 239 165 240
rect 165 239 166 240
rect 166 239 167 240
rect 167 239 168 240
rect 168 239 169 240
rect 169 239 170 240
rect 170 239 171 240
rect 171 239 172 240
rect 172 239 173 240
rect 173 239 174 240
rect 174 239 175 240
rect 175 239 176 240
rect 184 239 185 240
rect 185 239 186 240
rect 186 239 187 240
rect 187 239 188 240
rect 188 239 189 240
rect 189 239 190 240
rect 190 239 191 240
rect 193 239 194 240
rect 194 239 195 240
rect 195 239 196 240
rect 196 239 197 240
rect 197 239 198 240
rect 198 239 199 240
rect 199 239 200 240
rect 200 239 201 240
rect 201 239 202 240
rect 202 239 203 240
rect 203 239 204 240
rect 476 239 477 240
rect 477 239 478 240
rect 478 239 479 240
rect 479 239 480 240
rect 480 239 481 240
rect 481 239 482 240
rect 482 239 483 240
rect 483 239 484 240
rect 484 239 485 240
rect 485 239 486 240
rect 486 239 487 240
rect 487 239 488 240
rect 529 239 530 240
rect 530 239 531 240
rect 531 239 532 240
rect 532 239 533 240
rect 533 239 534 240
rect 534 239 535 240
rect 535 239 536 240
rect 536 239 537 240
rect 92 238 93 239
rect 93 238 94 239
rect 94 238 95 239
rect 95 238 96 239
rect 96 238 97 239
rect 118 238 119 239
rect 119 238 120 239
rect 120 238 121 239
rect 121 238 122 239
rect 122 238 123 239
rect 123 238 124 239
rect 124 238 125 239
rect 125 238 126 239
rect 126 238 127 239
rect 127 238 128 239
rect 128 238 129 239
rect 129 238 130 239
rect 130 238 131 239
rect 131 238 132 239
rect 132 238 133 239
rect 133 238 134 239
rect 134 238 135 239
rect 135 238 136 239
rect 136 238 137 239
rect 137 238 138 239
rect 138 238 139 239
rect 139 238 140 239
rect 140 238 141 239
rect 141 238 142 239
rect 142 238 143 239
rect 143 238 144 239
rect 154 238 155 239
rect 155 238 156 239
rect 156 238 157 239
rect 157 238 158 239
rect 158 238 159 239
rect 159 238 160 239
rect 160 238 161 239
rect 161 238 162 239
rect 162 238 163 239
rect 163 238 164 239
rect 164 238 165 239
rect 165 238 166 239
rect 166 238 167 239
rect 167 238 168 239
rect 168 238 169 239
rect 169 238 170 239
rect 170 238 171 239
rect 171 238 172 239
rect 172 238 173 239
rect 173 238 174 239
rect 174 238 175 239
rect 175 238 176 239
rect 176 238 177 239
rect 177 238 178 239
rect 178 238 179 239
rect 179 238 180 239
rect 180 238 181 239
rect 182 238 183 239
rect 183 238 184 239
rect 184 238 185 239
rect 185 238 186 239
rect 186 238 187 239
rect 187 238 188 239
rect 188 238 189 239
rect 189 238 190 239
rect 190 238 191 239
rect 193 238 194 239
rect 194 238 195 239
rect 195 238 196 239
rect 196 238 197 239
rect 197 238 198 239
rect 198 238 199 239
rect 199 238 200 239
rect 200 238 201 239
rect 201 238 202 239
rect 202 238 203 239
rect 203 238 204 239
rect 204 238 205 239
rect 205 238 206 239
rect 476 238 477 239
rect 477 238 478 239
rect 478 238 479 239
rect 479 238 480 239
rect 480 238 481 239
rect 481 238 482 239
rect 482 238 483 239
rect 483 238 484 239
rect 484 238 485 239
rect 485 238 486 239
rect 486 238 487 239
rect 487 238 488 239
rect 529 238 530 239
rect 530 238 531 239
rect 531 238 532 239
rect 532 238 533 239
rect 533 238 534 239
rect 534 238 535 239
rect 535 238 536 239
rect 536 238 537 239
rect 92 237 93 238
rect 93 237 94 238
rect 94 237 95 238
rect 95 237 96 238
rect 96 237 97 238
rect 118 237 119 238
rect 119 237 120 238
rect 120 237 121 238
rect 121 237 122 238
rect 122 237 123 238
rect 123 237 124 238
rect 124 237 125 238
rect 125 237 126 238
rect 126 237 127 238
rect 127 237 128 238
rect 128 237 129 238
rect 129 237 130 238
rect 130 237 131 238
rect 131 237 132 238
rect 132 237 133 238
rect 133 237 134 238
rect 134 237 135 238
rect 135 237 136 238
rect 136 237 137 238
rect 137 237 138 238
rect 138 237 139 238
rect 139 237 140 238
rect 140 237 141 238
rect 141 237 142 238
rect 142 237 143 238
rect 143 237 144 238
rect 154 237 155 238
rect 155 237 156 238
rect 156 237 157 238
rect 157 237 158 238
rect 158 237 159 238
rect 159 237 160 238
rect 160 237 161 238
rect 161 237 162 238
rect 162 237 163 238
rect 163 237 164 238
rect 164 237 165 238
rect 165 237 166 238
rect 166 237 167 238
rect 167 237 168 238
rect 168 237 169 238
rect 169 237 170 238
rect 170 237 171 238
rect 171 237 172 238
rect 172 237 173 238
rect 173 237 174 238
rect 174 237 175 238
rect 175 237 176 238
rect 176 237 177 238
rect 177 237 178 238
rect 178 237 179 238
rect 179 237 180 238
rect 180 237 181 238
rect 182 237 183 238
rect 183 237 184 238
rect 184 237 185 238
rect 185 237 186 238
rect 186 237 187 238
rect 187 237 188 238
rect 188 237 189 238
rect 193 237 194 238
rect 194 237 195 238
rect 195 237 196 238
rect 196 237 197 238
rect 197 237 198 238
rect 198 237 199 238
rect 199 237 200 238
rect 200 237 201 238
rect 201 237 202 238
rect 202 237 203 238
rect 203 237 204 238
rect 204 237 205 238
rect 205 237 206 238
rect 476 237 477 238
rect 477 237 478 238
rect 478 237 479 238
rect 479 237 480 238
rect 480 237 481 238
rect 481 237 482 238
rect 482 237 483 238
rect 483 237 484 238
rect 484 237 485 238
rect 485 237 486 238
rect 486 237 487 238
rect 487 237 488 238
rect 529 237 530 238
rect 530 237 531 238
rect 531 237 532 238
rect 532 237 533 238
rect 533 237 534 238
rect 534 237 535 238
rect 535 237 536 238
rect 536 237 537 238
rect 92 236 93 237
rect 93 236 94 237
rect 94 236 95 237
rect 95 236 96 237
rect 96 236 97 237
rect 118 236 119 237
rect 119 236 120 237
rect 120 236 121 237
rect 121 236 122 237
rect 122 236 123 237
rect 123 236 124 237
rect 124 236 125 237
rect 125 236 126 237
rect 126 236 127 237
rect 127 236 128 237
rect 128 236 129 237
rect 129 236 130 237
rect 130 236 131 237
rect 131 236 132 237
rect 132 236 133 237
rect 133 236 134 237
rect 134 236 135 237
rect 135 236 136 237
rect 136 236 137 237
rect 137 236 138 237
rect 138 236 139 237
rect 139 236 140 237
rect 140 236 141 237
rect 141 236 142 237
rect 142 236 143 237
rect 143 236 144 237
rect 152 236 153 237
rect 153 236 154 237
rect 154 236 155 237
rect 155 236 156 237
rect 156 236 157 237
rect 157 236 158 237
rect 158 236 159 237
rect 159 236 160 237
rect 160 236 161 237
rect 161 236 162 237
rect 162 236 163 237
rect 163 236 164 237
rect 164 236 165 237
rect 165 236 166 237
rect 166 236 167 237
rect 167 236 168 237
rect 168 236 169 237
rect 169 236 170 237
rect 170 236 171 237
rect 171 236 172 237
rect 172 236 173 237
rect 173 236 174 237
rect 174 236 175 237
rect 175 236 176 237
rect 176 236 177 237
rect 177 236 178 237
rect 178 236 179 237
rect 179 236 180 237
rect 180 236 181 237
rect 182 236 183 237
rect 183 236 184 237
rect 184 236 185 237
rect 185 236 186 237
rect 186 236 187 237
rect 187 236 188 237
rect 188 236 189 237
rect 193 236 194 237
rect 194 236 195 237
rect 195 236 196 237
rect 196 236 197 237
rect 197 236 198 237
rect 198 236 199 237
rect 199 236 200 237
rect 200 236 201 237
rect 201 236 202 237
rect 202 236 203 237
rect 203 236 204 237
rect 204 236 205 237
rect 205 236 206 237
rect 476 236 477 237
rect 477 236 478 237
rect 478 236 479 237
rect 479 236 480 237
rect 480 236 481 237
rect 481 236 482 237
rect 482 236 483 237
rect 483 236 484 237
rect 484 236 485 237
rect 485 236 486 237
rect 486 236 487 237
rect 487 236 488 237
rect 529 236 530 237
rect 530 236 531 237
rect 531 236 532 237
rect 532 236 533 237
rect 533 236 534 237
rect 534 236 535 237
rect 535 236 536 237
rect 536 236 537 237
rect 92 235 93 236
rect 93 235 94 236
rect 94 235 95 236
rect 95 235 96 236
rect 96 235 97 236
rect 120 235 121 236
rect 121 235 122 236
rect 122 235 123 236
rect 123 235 124 236
rect 124 235 125 236
rect 126 235 127 236
rect 127 235 128 236
rect 128 235 129 236
rect 129 235 130 236
rect 130 235 131 236
rect 132 235 133 236
rect 133 235 134 236
rect 134 235 135 236
rect 135 235 136 236
rect 137 235 138 236
rect 138 235 139 236
rect 139 235 140 236
rect 140 235 141 236
rect 141 235 142 236
rect 152 235 153 236
rect 153 235 154 236
rect 154 235 155 236
rect 156 235 157 236
rect 157 235 158 236
rect 158 235 159 236
rect 160 235 161 236
rect 161 235 162 236
rect 162 235 163 236
rect 163 235 164 236
rect 165 235 166 236
rect 166 235 167 236
rect 167 235 168 236
rect 168 235 169 236
rect 169 235 170 236
rect 171 235 172 236
rect 172 235 173 236
rect 173 235 174 236
rect 174 235 175 236
rect 175 235 176 236
rect 176 235 177 236
rect 177 235 178 236
rect 178 235 179 236
rect 179 235 180 236
rect 180 235 181 236
rect 182 235 183 236
rect 183 235 184 236
rect 184 235 185 236
rect 185 235 186 236
rect 186 235 187 236
rect 187 235 188 236
rect 188 235 189 236
rect 195 235 196 236
rect 196 235 197 236
rect 197 235 198 236
rect 198 235 199 236
rect 199 235 200 236
rect 200 235 201 236
rect 201 235 202 236
rect 202 235 203 236
rect 203 235 204 236
rect 204 235 205 236
rect 205 235 206 236
rect 476 235 477 236
rect 477 235 478 236
rect 478 235 479 236
rect 479 235 480 236
rect 480 235 481 236
rect 481 235 482 236
rect 482 235 483 236
rect 483 235 484 236
rect 484 235 485 236
rect 485 235 486 236
rect 486 235 487 236
rect 487 235 488 236
rect 529 235 530 236
rect 530 235 531 236
rect 531 235 532 236
rect 532 235 533 236
rect 533 235 534 236
rect 534 235 535 236
rect 535 235 536 236
rect 536 235 537 236
rect 92 234 93 235
rect 93 234 94 235
rect 94 234 95 235
rect 95 234 96 235
rect 96 234 97 235
rect 120 234 121 235
rect 121 234 122 235
rect 122 234 123 235
rect 123 234 124 235
rect 124 234 125 235
rect 126 234 127 235
rect 127 234 128 235
rect 128 234 129 235
rect 129 234 130 235
rect 130 234 131 235
rect 132 234 133 235
rect 133 234 134 235
rect 134 234 135 235
rect 135 234 136 235
rect 137 234 138 235
rect 138 234 139 235
rect 139 234 140 235
rect 140 234 141 235
rect 141 234 142 235
rect 152 234 153 235
rect 153 234 154 235
rect 154 234 155 235
rect 156 234 157 235
rect 157 234 158 235
rect 158 234 159 235
rect 160 234 161 235
rect 161 234 162 235
rect 162 234 163 235
rect 163 234 164 235
rect 165 234 166 235
rect 166 234 167 235
rect 167 234 168 235
rect 168 234 169 235
rect 169 234 170 235
rect 171 234 172 235
rect 172 234 173 235
rect 173 234 174 235
rect 174 234 175 235
rect 175 234 176 235
rect 176 234 177 235
rect 177 234 178 235
rect 178 234 179 235
rect 179 234 180 235
rect 180 234 181 235
rect 182 234 183 235
rect 183 234 184 235
rect 184 234 185 235
rect 185 234 186 235
rect 186 234 187 235
rect 187 234 188 235
rect 188 234 189 235
rect 195 234 196 235
rect 196 234 197 235
rect 197 234 198 235
rect 198 234 199 235
rect 199 234 200 235
rect 200 234 201 235
rect 201 234 202 235
rect 202 234 203 235
rect 203 234 204 235
rect 204 234 205 235
rect 205 234 206 235
rect 206 234 207 235
rect 414 234 415 235
rect 415 234 416 235
rect 416 234 417 235
rect 417 234 418 235
rect 418 234 419 235
rect 419 234 420 235
rect 420 234 421 235
rect 421 234 422 235
rect 422 234 423 235
rect 423 234 424 235
rect 424 234 425 235
rect 425 234 426 235
rect 426 234 427 235
rect 427 234 428 235
rect 428 234 429 235
rect 429 234 430 235
rect 430 234 431 235
rect 431 234 432 235
rect 432 234 433 235
rect 433 234 434 235
rect 434 234 435 235
rect 435 234 436 235
rect 436 234 437 235
rect 437 234 438 235
rect 438 234 439 235
rect 439 234 440 235
rect 440 234 441 235
rect 441 234 442 235
rect 442 234 443 235
rect 443 234 444 235
rect 444 234 445 235
rect 445 234 446 235
rect 446 234 447 235
rect 447 234 448 235
rect 448 234 449 235
rect 449 234 450 235
rect 450 234 451 235
rect 451 234 452 235
rect 452 234 453 235
rect 453 234 454 235
rect 454 234 455 235
rect 455 234 456 235
rect 456 234 457 235
rect 457 234 458 235
rect 458 234 459 235
rect 459 234 460 235
rect 460 234 461 235
rect 461 234 462 235
rect 462 234 463 235
rect 463 234 464 235
rect 464 234 465 235
rect 465 234 466 235
rect 476 234 477 235
rect 477 234 478 235
rect 478 234 479 235
rect 479 234 480 235
rect 480 234 481 235
rect 481 234 482 235
rect 482 234 483 235
rect 483 234 484 235
rect 484 234 485 235
rect 485 234 486 235
rect 486 234 487 235
rect 487 234 488 235
rect 527 234 528 235
rect 528 234 529 235
rect 529 234 530 235
rect 530 234 531 235
rect 531 234 532 235
rect 532 234 533 235
rect 533 234 534 235
rect 534 234 535 235
rect 535 234 536 235
rect 536 234 537 235
rect 92 233 93 234
rect 93 233 94 234
rect 94 233 95 234
rect 95 233 96 234
rect 96 233 97 234
rect 182 233 183 234
rect 183 233 184 234
rect 184 233 185 234
rect 185 233 186 234
rect 186 233 187 234
rect 195 233 196 234
rect 196 233 197 234
rect 197 233 198 234
rect 198 233 199 234
rect 199 233 200 234
rect 200 233 201 234
rect 201 233 202 234
rect 202 233 203 234
rect 203 233 204 234
rect 204 233 205 234
rect 205 233 206 234
rect 206 233 207 234
rect 414 233 415 234
rect 415 233 416 234
rect 416 233 417 234
rect 417 233 418 234
rect 418 233 419 234
rect 419 233 420 234
rect 420 233 421 234
rect 421 233 422 234
rect 422 233 423 234
rect 423 233 424 234
rect 424 233 425 234
rect 425 233 426 234
rect 426 233 427 234
rect 427 233 428 234
rect 428 233 429 234
rect 429 233 430 234
rect 430 233 431 234
rect 431 233 432 234
rect 432 233 433 234
rect 433 233 434 234
rect 434 233 435 234
rect 435 233 436 234
rect 436 233 437 234
rect 437 233 438 234
rect 438 233 439 234
rect 439 233 440 234
rect 440 233 441 234
rect 441 233 442 234
rect 442 233 443 234
rect 443 233 444 234
rect 444 233 445 234
rect 445 233 446 234
rect 446 233 447 234
rect 447 233 448 234
rect 448 233 449 234
rect 449 233 450 234
rect 450 233 451 234
rect 451 233 452 234
rect 452 233 453 234
rect 453 233 454 234
rect 454 233 455 234
rect 455 233 456 234
rect 456 233 457 234
rect 457 233 458 234
rect 458 233 459 234
rect 459 233 460 234
rect 460 233 461 234
rect 461 233 462 234
rect 462 233 463 234
rect 463 233 464 234
rect 464 233 465 234
rect 465 233 466 234
rect 476 233 477 234
rect 477 233 478 234
rect 478 233 479 234
rect 479 233 480 234
rect 480 233 481 234
rect 481 233 482 234
rect 482 233 483 234
rect 483 233 484 234
rect 484 233 485 234
rect 485 233 486 234
rect 486 233 487 234
rect 487 233 488 234
rect 527 233 528 234
rect 528 233 529 234
rect 529 233 530 234
rect 530 233 531 234
rect 531 233 532 234
rect 532 233 533 234
rect 533 233 534 234
rect 534 233 535 234
rect 535 233 536 234
rect 536 233 537 234
rect 92 232 93 233
rect 93 232 94 233
rect 94 232 95 233
rect 95 232 96 233
rect 96 232 97 233
rect 180 232 181 233
rect 181 232 182 233
rect 182 232 183 233
rect 183 232 184 233
rect 184 232 185 233
rect 185 232 186 233
rect 186 232 187 233
rect 195 232 196 233
rect 196 232 197 233
rect 197 232 198 233
rect 198 232 199 233
rect 199 232 200 233
rect 200 232 201 233
rect 201 232 202 233
rect 202 232 203 233
rect 203 232 204 233
rect 204 232 205 233
rect 205 232 206 233
rect 206 232 207 233
rect 414 232 415 233
rect 415 232 416 233
rect 416 232 417 233
rect 417 232 418 233
rect 418 232 419 233
rect 419 232 420 233
rect 420 232 421 233
rect 421 232 422 233
rect 422 232 423 233
rect 423 232 424 233
rect 424 232 425 233
rect 425 232 426 233
rect 426 232 427 233
rect 427 232 428 233
rect 428 232 429 233
rect 429 232 430 233
rect 430 232 431 233
rect 431 232 432 233
rect 432 232 433 233
rect 433 232 434 233
rect 434 232 435 233
rect 435 232 436 233
rect 436 232 437 233
rect 437 232 438 233
rect 438 232 439 233
rect 439 232 440 233
rect 440 232 441 233
rect 441 232 442 233
rect 442 232 443 233
rect 443 232 444 233
rect 444 232 445 233
rect 445 232 446 233
rect 446 232 447 233
rect 447 232 448 233
rect 448 232 449 233
rect 449 232 450 233
rect 450 232 451 233
rect 451 232 452 233
rect 452 232 453 233
rect 453 232 454 233
rect 454 232 455 233
rect 455 232 456 233
rect 456 232 457 233
rect 457 232 458 233
rect 458 232 459 233
rect 459 232 460 233
rect 460 232 461 233
rect 461 232 462 233
rect 462 232 463 233
rect 463 232 464 233
rect 464 232 465 233
rect 465 232 466 233
rect 466 232 467 233
rect 467 232 468 233
rect 476 232 477 233
rect 477 232 478 233
rect 478 232 479 233
rect 479 232 480 233
rect 480 232 481 233
rect 481 232 482 233
rect 482 232 483 233
rect 483 232 484 233
rect 484 232 485 233
rect 485 232 486 233
rect 486 232 487 233
rect 487 232 488 233
rect 527 232 528 233
rect 528 232 529 233
rect 529 232 530 233
rect 530 232 531 233
rect 531 232 532 233
rect 532 232 533 233
rect 533 232 534 233
rect 534 232 535 233
rect 535 232 536 233
rect 536 232 537 233
rect 92 231 93 232
rect 93 231 94 232
rect 94 231 95 232
rect 95 231 96 232
rect 96 231 97 232
rect 180 231 181 232
rect 181 231 182 232
rect 182 231 183 232
rect 183 231 184 232
rect 184 231 185 232
rect 185 231 186 232
rect 186 231 187 232
rect 197 231 198 232
rect 198 231 199 232
rect 199 231 200 232
rect 200 231 201 232
rect 201 231 202 232
rect 202 231 203 232
rect 203 231 204 232
rect 204 231 205 232
rect 205 231 206 232
rect 206 231 207 232
rect 414 231 415 232
rect 415 231 416 232
rect 416 231 417 232
rect 417 231 418 232
rect 418 231 419 232
rect 419 231 420 232
rect 420 231 421 232
rect 421 231 422 232
rect 422 231 423 232
rect 423 231 424 232
rect 424 231 425 232
rect 425 231 426 232
rect 426 231 427 232
rect 427 231 428 232
rect 428 231 429 232
rect 429 231 430 232
rect 430 231 431 232
rect 431 231 432 232
rect 432 231 433 232
rect 433 231 434 232
rect 434 231 435 232
rect 435 231 436 232
rect 436 231 437 232
rect 437 231 438 232
rect 438 231 439 232
rect 439 231 440 232
rect 440 231 441 232
rect 441 231 442 232
rect 442 231 443 232
rect 443 231 444 232
rect 444 231 445 232
rect 445 231 446 232
rect 446 231 447 232
rect 447 231 448 232
rect 448 231 449 232
rect 449 231 450 232
rect 450 231 451 232
rect 451 231 452 232
rect 452 231 453 232
rect 453 231 454 232
rect 454 231 455 232
rect 455 231 456 232
rect 456 231 457 232
rect 457 231 458 232
rect 458 231 459 232
rect 459 231 460 232
rect 460 231 461 232
rect 461 231 462 232
rect 462 231 463 232
rect 463 231 464 232
rect 464 231 465 232
rect 465 231 466 232
rect 466 231 467 232
rect 467 231 468 232
rect 476 231 477 232
rect 477 231 478 232
rect 478 231 479 232
rect 479 231 480 232
rect 480 231 481 232
rect 481 231 482 232
rect 482 231 483 232
rect 483 231 484 232
rect 484 231 485 232
rect 485 231 486 232
rect 486 231 487 232
rect 527 231 528 232
rect 528 231 529 232
rect 529 231 530 232
rect 530 231 531 232
rect 531 231 532 232
rect 532 231 533 232
rect 533 231 534 232
rect 534 231 535 232
rect 92 230 93 231
rect 93 230 94 231
rect 94 230 95 231
rect 95 230 96 231
rect 96 230 97 231
rect 180 230 181 231
rect 181 230 182 231
rect 182 230 183 231
rect 183 230 184 231
rect 184 230 185 231
rect 185 230 186 231
rect 186 230 187 231
rect 197 230 198 231
rect 198 230 199 231
rect 199 230 200 231
rect 200 230 201 231
rect 201 230 202 231
rect 202 230 203 231
rect 203 230 204 231
rect 204 230 205 231
rect 205 230 206 231
rect 206 230 207 231
rect 414 230 415 231
rect 415 230 416 231
rect 416 230 417 231
rect 417 230 418 231
rect 418 230 419 231
rect 419 230 420 231
rect 420 230 421 231
rect 421 230 422 231
rect 422 230 423 231
rect 423 230 424 231
rect 424 230 425 231
rect 425 230 426 231
rect 426 230 427 231
rect 427 230 428 231
rect 428 230 429 231
rect 429 230 430 231
rect 430 230 431 231
rect 431 230 432 231
rect 432 230 433 231
rect 433 230 434 231
rect 434 230 435 231
rect 435 230 436 231
rect 436 230 437 231
rect 437 230 438 231
rect 438 230 439 231
rect 439 230 440 231
rect 440 230 441 231
rect 441 230 442 231
rect 442 230 443 231
rect 443 230 444 231
rect 444 230 445 231
rect 445 230 446 231
rect 446 230 447 231
rect 447 230 448 231
rect 448 230 449 231
rect 449 230 450 231
rect 450 230 451 231
rect 451 230 452 231
rect 452 230 453 231
rect 453 230 454 231
rect 454 230 455 231
rect 455 230 456 231
rect 456 230 457 231
rect 457 230 458 231
rect 458 230 459 231
rect 459 230 460 231
rect 460 230 461 231
rect 461 230 462 231
rect 462 230 463 231
rect 463 230 464 231
rect 464 230 465 231
rect 465 230 466 231
rect 466 230 467 231
rect 467 230 468 231
rect 476 230 477 231
rect 477 230 478 231
rect 478 230 479 231
rect 479 230 480 231
rect 480 230 481 231
rect 481 230 482 231
rect 482 230 483 231
rect 483 230 484 231
rect 484 230 485 231
rect 485 230 486 231
rect 486 230 487 231
rect 527 230 528 231
rect 528 230 529 231
rect 529 230 530 231
rect 530 230 531 231
rect 531 230 532 231
rect 532 230 533 231
rect 533 230 534 231
rect 534 230 535 231
rect 90 229 91 230
rect 91 229 92 230
rect 92 229 93 230
rect 93 229 94 230
rect 94 229 95 230
rect 95 229 96 230
rect 96 229 97 230
rect 180 229 181 230
rect 181 229 182 230
rect 182 229 183 230
rect 183 229 184 230
rect 184 229 185 230
rect 185 229 186 230
rect 186 229 187 230
rect 197 229 198 230
rect 198 229 199 230
rect 199 229 200 230
rect 200 229 201 230
rect 201 229 202 230
rect 202 229 203 230
rect 203 229 204 230
rect 204 229 205 230
rect 205 229 206 230
rect 206 229 207 230
rect 207 229 208 230
rect 208 229 209 230
rect 414 229 415 230
rect 415 229 416 230
rect 416 229 417 230
rect 417 229 418 230
rect 418 229 419 230
rect 419 229 420 230
rect 420 229 421 230
rect 421 229 422 230
rect 422 229 423 230
rect 423 229 424 230
rect 424 229 425 230
rect 425 229 426 230
rect 426 229 427 230
rect 427 229 428 230
rect 428 229 429 230
rect 429 229 430 230
rect 430 229 431 230
rect 431 229 432 230
rect 432 229 433 230
rect 433 229 434 230
rect 434 229 435 230
rect 435 229 436 230
rect 436 229 437 230
rect 437 229 438 230
rect 438 229 439 230
rect 439 229 440 230
rect 440 229 441 230
rect 441 229 442 230
rect 442 229 443 230
rect 443 229 444 230
rect 444 229 445 230
rect 445 229 446 230
rect 446 229 447 230
rect 447 229 448 230
rect 448 229 449 230
rect 449 229 450 230
rect 450 229 451 230
rect 451 229 452 230
rect 452 229 453 230
rect 453 229 454 230
rect 454 229 455 230
rect 455 229 456 230
rect 456 229 457 230
rect 457 229 458 230
rect 458 229 459 230
rect 459 229 460 230
rect 460 229 461 230
rect 461 229 462 230
rect 462 229 463 230
rect 463 229 464 230
rect 464 229 465 230
rect 465 229 466 230
rect 466 229 467 230
rect 467 229 468 230
rect 476 229 477 230
rect 477 229 478 230
rect 478 229 479 230
rect 479 229 480 230
rect 480 229 481 230
rect 481 229 482 230
rect 482 229 483 230
rect 483 229 484 230
rect 484 229 485 230
rect 485 229 486 230
rect 486 229 487 230
rect 487 229 488 230
rect 527 229 528 230
rect 528 229 529 230
rect 529 229 530 230
rect 530 229 531 230
rect 531 229 532 230
rect 532 229 533 230
rect 533 229 534 230
rect 534 229 535 230
rect 90 228 91 229
rect 91 228 92 229
rect 92 228 93 229
rect 93 228 94 229
rect 94 228 95 229
rect 95 228 96 229
rect 96 228 97 229
rect 180 228 181 229
rect 181 228 182 229
rect 182 228 183 229
rect 183 228 184 229
rect 184 228 185 229
rect 185 228 186 229
rect 186 228 187 229
rect 197 228 198 229
rect 198 228 199 229
rect 199 228 200 229
rect 200 228 201 229
rect 201 228 202 229
rect 202 228 203 229
rect 203 228 204 229
rect 204 228 205 229
rect 205 228 206 229
rect 206 228 207 229
rect 207 228 208 229
rect 208 228 209 229
rect 414 228 415 229
rect 415 228 416 229
rect 416 228 417 229
rect 417 228 418 229
rect 418 228 419 229
rect 419 228 420 229
rect 420 228 421 229
rect 421 228 422 229
rect 422 228 423 229
rect 423 228 424 229
rect 424 228 425 229
rect 425 228 426 229
rect 426 228 427 229
rect 427 228 428 229
rect 429 228 430 229
rect 430 228 431 229
rect 431 228 432 229
rect 433 228 434 229
rect 434 228 435 229
rect 435 228 436 229
rect 436 228 437 229
rect 437 228 438 229
rect 438 228 439 229
rect 439 228 440 229
rect 440 228 441 229
rect 441 228 442 229
rect 442 228 443 229
rect 443 228 444 229
rect 444 228 445 229
rect 446 228 447 229
rect 447 228 448 229
rect 448 228 449 229
rect 449 228 450 229
rect 450 228 451 229
rect 452 228 453 229
rect 453 228 454 229
rect 454 228 455 229
rect 455 228 456 229
rect 456 228 457 229
rect 457 228 458 229
rect 458 228 459 229
rect 459 228 460 229
rect 460 228 461 229
rect 461 228 462 229
rect 462 228 463 229
rect 463 228 464 229
rect 464 228 465 229
rect 465 228 466 229
rect 476 228 477 229
rect 477 228 478 229
rect 478 228 479 229
rect 479 228 480 229
rect 480 228 481 229
rect 481 228 482 229
rect 482 228 483 229
rect 483 228 484 229
rect 484 228 485 229
rect 485 228 486 229
rect 486 228 487 229
rect 487 228 488 229
rect 527 228 528 229
rect 528 228 529 229
rect 529 228 530 229
rect 530 228 531 229
rect 531 228 532 229
rect 532 228 533 229
rect 533 228 534 229
rect 534 228 535 229
rect 90 227 91 228
rect 91 227 92 228
rect 92 227 93 228
rect 93 227 94 228
rect 94 227 95 228
rect 95 227 96 228
rect 96 227 97 228
rect 178 227 179 228
rect 179 227 180 228
rect 180 227 181 228
rect 181 227 182 228
rect 182 227 183 228
rect 183 227 184 228
rect 184 227 185 228
rect 185 227 186 228
rect 186 227 187 228
rect 197 227 198 228
rect 198 227 199 228
rect 199 227 200 228
rect 200 227 201 228
rect 201 227 202 228
rect 202 227 203 228
rect 203 227 204 228
rect 204 227 205 228
rect 205 227 206 228
rect 206 227 207 228
rect 207 227 208 228
rect 208 227 209 228
rect 414 227 415 228
rect 415 227 416 228
rect 416 227 417 228
rect 417 227 418 228
rect 418 227 419 228
rect 419 227 420 228
rect 420 227 421 228
rect 421 227 422 228
rect 422 227 423 228
rect 423 227 424 228
rect 424 227 425 228
rect 425 227 426 228
rect 426 227 427 228
rect 427 227 428 228
rect 429 227 430 228
rect 430 227 431 228
rect 431 227 432 228
rect 433 227 434 228
rect 434 227 435 228
rect 435 227 436 228
rect 436 227 437 228
rect 437 227 438 228
rect 438 227 439 228
rect 439 227 440 228
rect 440 227 441 228
rect 441 227 442 228
rect 442 227 443 228
rect 443 227 444 228
rect 444 227 445 228
rect 446 227 447 228
rect 447 227 448 228
rect 448 227 449 228
rect 449 227 450 228
rect 450 227 451 228
rect 452 227 453 228
rect 453 227 454 228
rect 454 227 455 228
rect 455 227 456 228
rect 456 227 457 228
rect 457 227 458 228
rect 458 227 459 228
rect 459 227 460 228
rect 460 227 461 228
rect 461 227 462 228
rect 462 227 463 228
rect 463 227 464 228
rect 464 227 465 228
rect 465 227 466 228
rect 476 227 477 228
rect 477 227 478 228
rect 478 227 479 228
rect 479 227 480 228
rect 480 227 481 228
rect 481 227 482 228
rect 482 227 483 228
rect 483 227 484 228
rect 484 227 485 228
rect 485 227 486 228
rect 486 227 487 228
rect 487 227 488 228
rect 527 227 528 228
rect 528 227 529 228
rect 529 227 530 228
rect 530 227 531 228
rect 531 227 532 228
rect 532 227 533 228
rect 533 227 534 228
rect 534 227 535 228
rect 90 226 91 227
rect 91 226 92 227
rect 92 226 93 227
rect 93 226 94 227
rect 94 226 95 227
rect 95 226 96 227
rect 96 226 97 227
rect 178 226 179 227
rect 179 226 180 227
rect 180 226 181 227
rect 181 226 182 227
rect 182 226 183 227
rect 183 226 184 227
rect 184 226 185 227
rect 199 226 200 227
rect 200 226 201 227
rect 201 226 202 227
rect 202 226 203 227
rect 203 226 204 227
rect 204 226 205 227
rect 205 226 206 227
rect 206 226 207 227
rect 207 226 208 227
rect 208 226 209 227
rect 414 226 415 227
rect 415 226 416 227
rect 416 226 417 227
rect 417 226 418 227
rect 418 226 419 227
rect 419 226 420 227
rect 420 226 421 227
rect 421 226 422 227
rect 422 226 423 227
rect 435 226 436 227
rect 436 226 437 227
rect 437 226 438 227
rect 438 226 439 227
rect 439 226 440 227
rect 440 226 441 227
rect 441 226 442 227
rect 442 226 443 227
rect 443 226 444 227
rect 444 226 445 227
rect 457 226 458 227
rect 458 226 459 227
rect 459 226 460 227
rect 460 226 461 227
rect 461 226 462 227
rect 462 226 463 227
rect 463 226 464 227
rect 464 226 465 227
rect 465 226 466 227
rect 476 226 477 227
rect 477 226 478 227
rect 478 226 479 227
rect 479 226 480 227
rect 480 226 481 227
rect 481 226 482 227
rect 482 226 483 227
rect 483 226 484 227
rect 484 226 485 227
rect 485 226 486 227
rect 486 226 487 227
rect 487 226 488 227
rect 527 226 528 227
rect 528 226 529 227
rect 529 226 530 227
rect 530 226 531 227
rect 531 226 532 227
rect 532 226 533 227
rect 533 226 534 227
rect 534 226 535 227
rect 88 225 89 226
rect 89 225 90 226
rect 90 225 91 226
rect 91 225 92 226
rect 92 225 93 226
rect 93 225 94 226
rect 94 225 95 226
rect 95 225 96 226
rect 96 225 97 226
rect 97 225 98 226
rect 98 225 99 226
rect 178 225 179 226
rect 179 225 180 226
rect 180 225 181 226
rect 181 225 182 226
rect 182 225 183 226
rect 183 225 184 226
rect 184 225 185 226
rect 199 225 200 226
rect 200 225 201 226
rect 201 225 202 226
rect 202 225 203 226
rect 203 225 204 226
rect 204 225 205 226
rect 205 225 206 226
rect 206 225 207 226
rect 207 225 208 226
rect 208 225 209 226
rect 414 225 415 226
rect 415 225 416 226
rect 416 225 417 226
rect 417 225 418 226
rect 418 225 419 226
rect 419 225 420 226
rect 420 225 421 226
rect 421 225 422 226
rect 422 225 423 226
rect 435 225 436 226
rect 436 225 437 226
rect 437 225 438 226
rect 438 225 439 226
rect 439 225 440 226
rect 440 225 441 226
rect 441 225 442 226
rect 442 225 443 226
rect 443 225 444 226
rect 444 225 445 226
rect 457 225 458 226
rect 458 225 459 226
rect 459 225 460 226
rect 460 225 461 226
rect 461 225 462 226
rect 462 225 463 226
rect 463 225 464 226
rect 464 225 465 226
rect 465 225 466 226
rect 476 225 477 226
rect 477 225 478 226
rect 478 225 479 226
rect 479 225 480 226
rect 480 225 481 226
rect 481 225 482 226
rect 482 225 483 226
rect 483 225 484 226
rect 484 225 485 226
rect 485 225 486 226
rect 486 225 487 226
rect 487 225 488 226
rect 525 225 526 226
rect 526 225 527 226
rect 527 225 528 226
rect 528 225 529 226
rect 529 225 530 226
rect 530 225 531 226
rect 531 225 532 226
rect 532 225 533 226
rect 533 225 534 226
rect 534 225 535 226
rect 88 224 89 225
rect 89 224 90 225
rect 90 224 91 225
rect 91 224 92 225
rect 92 224 93 225
rect 93 224 94 225
rect 94 224 95 225
rect 95 224 96 225
rect 96 224 97 225
rect 97 224 98 225
rect 98 224 99 225
rect 178 224 179 225
rect 179 224 180 225
rect 180 224 181 225
rect 181 224 182 225
rect 182 224 183 225
rect 183 224 184 225
rect 184 224 185 225
rect 199 224 200 225
rect 200 224 201 225
rect 201 224 202 225
rect 202 224 203 225
rect 203 224 204 225
rect 204 224 205 225
rect 205 224 206 225
rect 206 224 207 225
rect 207 224 208 225
rect 208 224 209 225
rect 414 224 415 225
rect 415 224 416 225
rect 416 224 417 225
rect 417 224 418 225
rect 418 224 419 225
rect 419 224 420 225
rect 420 224 421 225
rect 435 224 436 225
rect 436 224 437 225
rect 437 224 438 225
rect 438 224 439 225
rect 439 224 440 225
rect 440 224 441 225
rect 441 224 442 225
rect 442 224 443 225
rect 443 224 444 225
rect 444 224 445 225
rect 461 224 462 225
rect 462 224 463 225
rect 463 224 464 225
rect 464 224 465 225
rect 465 224 466 225
rect 476 224 477 225
rect 477 224 478 225
rect 478 224 479 225
rect 479 224 480 225
rect 480 224 481 225
rect 481 224 482 225
rect 482 224 483 225
rect 483 224 484 225
rect 484 224 485 225
rect 485 224 486 225
rect 486 224 487 225
rect 525 224 526 225
rect 526 224 527 225
rect 527 224 528 225
rect 528 224 529 225
rect 529 224 530 225
rect 530 224 531 225
rect 531 224 532 225
rect 532 224 533 225
rect 533 224 534 225
rect 534 224 535 225
rect 88 223 89 224
rect 89 223 90 224
rect 90 223 91 224
rect 91 223 92 224
rect 92 223 93 224
rect 93 223 94 224
rect 94 223 95 224
rect 95 223 96 224
rect 96 223 97 224
rect 97 223 98 224
rect 98 223 99 224
rect 178 223 179 224
rect 179 223 180 224
rect 180 223 181 224
rect 181 223 182 224
rect 182 223 183 224
rect 183 223 184 224
rect 184 223 185 224
rect 199 223 200 224
rect 200 223 201 224
rect 201 223 202 224
rect 202 223 203 224
rect 203 223 204 224
rect 204 223 205 224
rect 205 223 206 224
rect 206 223 207 224
rect 207 223 208 224
rect 208 223 209 224
rect 209 223 210 224
rect 210 223 211 224
rect 412 223 413 224
rect 413 223 414 224
rect 414 223 415 224
rect 415 223 416 224
rect 416 223 417 224
rect 417 223 418 224
rect 418 223 419 224
rect 419 223 420 224
rect 420 223 421 224
rect 433 223 434 224
rect 434 223 435 224
rect 435 223 436 224
rect 436 223 437 224
rect 437 223 438 224
rect 438 223 439 224
rect 439 223 440 224
rect 440 223 441 224
rect 441 223 442 224
rect 442 223 443 224
rect 443 223 444 224
rect 444 223 445 224
rect 461 223 462 224
rect 462 223 463 224
rect 463 223 464 224
rect 464 223 465 224
rect 465 223 466 224
rect 476 223 477 224
rect 477 223 478 224
rect 478 223 479 224
rect 479 223 480 224
rect 480 223 481 224
rect 481 223 482 224
rect 482 223 483 224
rect 483 223 484 224
rect 484 223 485 224
rect 485 223 486 224
rect 486 223 487 224
rect 487 223 488 224
rect 525 223 526 224
rect 526 223 527 224
rect 527 223 528 224
rect 528 223 529 224
rect 529 223 530 224
rect 530 223 531 224
rect 531 223 532 224
rect 532 223 533 224
rect 533 223 534 224
rect 534 223 535 224
rect 90 222 91 223
rect 91 222 92 223
rect 92 222 93 223
rect 93 222 94 223
rect 94 222 95 223
rect 95 222 96 223
rect 96 222 97 223
rect 97 222 98 223
rect 98 222 99 223
rect 178 222 179 223
rect 179 222 180 223
rect 180 222 181 223
rect 181 222 182 223
rect 182 222 183 223
rect 199 222 200 223
rect 200 222 201 223
rect 201 222 202 223
rect 202 222 203 223
rect 203 222 204 223
rect 204 222 205 223
rect 205 222 206 223
rect 206 222 207 223
rect 207 222 208 223
rect 208 222 209 223
rect 209 222 210 223
rect 210 222 211 223
rect 412 222 413 223
rect 413 222 414 223
rect 414 222 415 223
rect 415 222 416 223
rect 416 222 417 223
rect 417 222 418 223
rect 418 222 419 223
rect 433 222 434 223
rect 434 222 435 223
rect 435 222 436 223
rect 436 222 437 223
rect 437 222 438 223
rect 438 222 439 223
rect 439 222 440 223
rect 440 222 441 223
rect 441 222 442 223
rect 442 222 443 223
rect 443 222 444 223
rect 444 222 445 223
rect 461 222 462 223
rect 462 222 463 223
rect 463 222 464 223
rect 464 222 465 223
rect 465 222 466 223
rect 476 222 477 223
rect 477 222 478 223
rect 478 222 479 223
rect 479 222 480 223
rect 480 222 481 223
rect 481 222 482 223
rect 482 222 483 223
rect 483 222 484 223
rect 484 222 485 223
rect 485 222 486 223
rect 486 222 487 223
rect 487 222 488 223
rect 525 222 526 223
rect 526 222 527 223
rect 527 222 528 223
rect 528 222 529 223
rect 529 222 530 223
rect 530 222 531 223
rect 531 222 532 223
rect 532 222 533 223
rect 533 222 534 223
rect 534 222 535 223
rect 90 221 91 222
rect 91 221 92 222
rect 92 221 93 222
rect 93 221 94 222
rect 94 221 95 222
rect 95 221 96 222
rect 96 221 97 222
rect 97 221 98 222
rect 98 221 99 222
rect 176 221 177 222
rect 177 221 178 222
rect 178 221 179 222
rect 179 221 180 222
rect 180 221 181 222
rect 181 221 182 222
rect 182 221 183 222
rect 183 221 184 222
rect 184 221 185 222
rect 185 221 186 222
rect 186 221 187 222
rect 190 221 191 222
rect 191 221 192 222
rect 195 221 196 222
rect 196 221 197 222
rect 197 221 198 222
rect 199 221 200 222
rect 200 221 201 222
rect 201 221 202 222
rect 202 221 203 222
rect 203 221 204 222
rect 204 221 205 222
rect 205 221 206 222
rect 206 221 207 222
rect 207 221 208 222
rect 208 221 209 222
rect 209 221 210 222
rect 210 221 211 222
rect 412 221 413 222
rect 413 221 414 222
rect 414 221 415 222
rect 415 221 416 222
rect 416 221 417 222
rect 417 221 418 222
rect 418 221 419 222
rect 433 221 434 222
rect 434 221 435 222
rect 435 221 436 222
rect 436 221 437 222
rect 437 221 438 222
rect 438 221 439 222
rect 439 221 440 222
rect 440 221 441 222
rect 441 221 442 222
rect 442 221 443 222
rect 443 221 444 222
rect 444 221 445 222
rect 461 221 462 222
rect 462 221 463 222
rect 463 221 464 222
rect 464 221 465 222
rect 465 221 466 222
rect 466 221 467 222
rect 467 221 468 222
rect 476 221 477 222
rect 477 221 478 222
rect 478 221 479 222
rect 479 221 480 222
rect 480 221 481 222
rect 481 221 482 222
rect 482 221 483 222
rect 483 221 484 222
rect 484 221 485 222
rect 485 221 486 222
rect 486 221 487 222
rect 487 221 488 222
rect 525 221 526 222
rect 526 221 527 222
rect 527 221 528 222
rect 528 221 529 222
rect 529 221 530 222
rect 530 221 531 222
rect 531 221 532 222
rect 532 221 533 222
rect 533 221 534 222
rect 534 221 535 222
rect 90 220 91 221
rect 91 220 92 221
rect 92 220 93 221
rect 93 220 94 221
rect 94 220 95 221
rect 95 220 96 221
rect 96 220 97 221
rect 97 220 98 221
rect 98 220 99 221
rect 176 220 177 221
rect 177 220 178 221
rect 178 220 179 221
rect 179 220 180 221
rect 180 220 181 221
rect 181 220 182 221
rect 182 220 183 221
rect 183 220 184 221
rect 184 220 185 221
rect 185 220 186 221
rect 186 220 187 221
rect 190 220 191 221
rect 191 220 192 221
rect 195 220 196 221
rect 196 220 197 221
rect 197 220 198 221
rect 201 220 202 221
rect 202 220 203 221
rect 203 220 204 221
rect 204 220 205 221
rect 205 220 206 221
rect 206 220 207 221
rect 207 220 208 221
rect 208 220 209 221
rect 209 220 210 221
rect 210 220 211 221
rect 414 220 415 221
rect 415 220 416 221
rect 416 220 417 221
rect 417 220 418 221
rect 418 220 419 221
rect 435 220 436 221
rect 436 220 437 221
rect 437 220 438 221
rect 438 220 439 221
rect 439 220 440 221
rect 440 220 441 221
rect 441 220 442 221
rect 442 220 443 221
rect 443 220 444 221
rect 444 220 445 221
rect 461 220 462 221
rect 462 220 463 221
rect 463 220 464 221
rect 464 220 465 221
rect 465 220 466 221
rect 466 220 467 221
rect 467 220 468 221
rect 476 220 477 221
rect 477 220 478 221
rect 478 220 479 221
rect 479 220 480 221
rect 480 220 481 221
rect 481 220 482 221
rect 482 220 483 221
rect 483 220 484 221
rect 484 220 485 221
rect 485 220 486 221
rect 486 220 487 221
rect 487 220 488 221
rect 525 220 526 221
rect 526 220 527 221
rect 527 220 528 221
rect 528 220 529 221
rect 529 220 530 221
rect 530 220 531 221
rect 531 220 532 221
rect 532 220 533 221
rect 90 219 91 220
rect 91 219 92 220
rect 92 219 93 220
rect 93 219 94 220
rect 94 219 95 220
rect 95 219 96 220
rect 96 219 97 220
rect 97 219 98 220
rect 98 219 99 220
rect 176 219 177 220
rect 177 219 178 220
rect 178 219 179 220
rect 179 219 180 220
rect 180 219 181 220
rect 181 219 182 220
rect 182 219 183 220
rect 183 219 184 220
rect 184 219 185 220
rect 185 219 186 220
rect 186 219 187 220
rect 187 219 188 220
rect 188 219 189 220
rect 189 219 190 220
rect 190 219 191 220
rect 191 219 192 220
rect 192 219 193 220
rect 193 219 194 220
rect 194 219 195 220
rect 195 219 196 220
rect 196 219 197 220
rect 197 219 198 220
rect 198 219 199 220
rect 199 219 200 220
rect 200 219 201 220
rect 201 219 202 220
rect 202 219 203 220
rect 203 219 204 220
rect 204 219 205 220
rect 205 219 206 220
rect 206 219 207 220
rect 207 219 208 220
rect 208 219 209 220
rect 209 219 210 220
rect 210 219 211 220
rect 211 219 212 220
rect 212 219 213 220
rect 414 219 415 220
rect 415 219 416 220
rect 416 219 417 220
rect 417 219 418 220
rect 418 219 419 220
rect 435 219 436 220
rect 436 219 437 220
rect 437 219 438 220
rect 438 219 439 220
rect 439 219 440 220
rect 440 219 441 220
rect 441 219 442 220
rect 442 219 443 220
rect 443 219 444 220
rect 444 219 445 220
rect 461 219 462 220
rect 462 219 463 220
rect 463 219 464 220
rect 464 219 465 220
rect 465 219 466 220
rect 466 219 467 220
rect 467 219 468 220
rect 476 219 477 220
rect 477 219 478 220
rect 478 219 479 220
rect 479 219 480 220
rect 480 219 481 220
rect 481 219 482 220
rect 482 219 483 220
rect 483 219 484 220
rect 484 219 485 220
rect 485 219 486 220
rect 486 219 487 220
rect 487 219 488 220
rect 523 219 524 220
rect 524 219 525 220
rect 525 219 526 220
rect 526 219 527 220
rect 527 219 528 220
rect 528 219 529 220
rect 529 219 530 220
rect 530 219 531 220
rect 531 219 532 220
rect 532 219 533 220
rect 90 218 91 219
rect 91 218 92 219
rect 92 218 93 219
rect 93 218 94 219
rect 94 218 95 219
rect 95 218 96 219
rect 96 218 97 219
rect 97 218 98 219
rect 98 218 99 219
rect 176 218 177 219
rect 177 218 178 219
rect 178 218 179 219
rect 179 218 180 219
rect 180 218 181 219
rect 181 218 182 219
rect 182 218 183 219
rect 183 218 184 219
rect 184 218 185 219
rect 185 218 186 219
rect 186 218 187 219
rect 187 218 188 219
rect 188 218 189 219
rect 189 218 190 219
rect 190 218 191 219
rect 191 218 192 219
rect 192 218 193 219
rect 193 218 194 219
rect 194 218 195 219
rect 195 218 196 219
rect 196 218 197 219
rect 197 218 198 219
rect 198 218 199 219
rect 199 218 200 219
rect 200 218 201 219
rect 201 218 202 219
rect 202 218 203 219
rect 203 218 204 219
rect 204 218 205 219
rect 205 218 206 219
rect 206 218 207 219
rect 207 218 208 219
rect 208 218 209 219
rect 209 218 210 219
rect 210 218 211 219
rect 211 218 212 219
rect 212 218 213 219
rect 414 218 415 219
rect 415 218 416 219
rect 416 218 417 219
rect 435 218 436 219
rect 436 218 437 219
rect 437 218 438 219
rect 438 218 439 219
rect 439 218 440 219
rect 440 218 441 219
rect 441 218 442 219
rect 442 218 443 219
rect 443 218 444 219
rect 444 218 445 219
rect 461 218 462 219
rect 462 218 463 219
rect 463 218 464 219
rect 464 218 465 219
rect 465 218 466 219
rect 476 218 477 219
rect 477 218 478 219
rect 478 218 479 219
rect 479 218 480 219
rect 480 218 481 219
rect 481 218 482 219
rect 482 218 483 219
rect 483 218 484 219
rect 484 218 485 219
rect 485 218 486 219
rect 486 218 487 219
rect 487 218 488 219
rect 523 218 524 219
rect 524 218 525 219
rect 525 218 526 219
rect 526 218 527 219
rect 527 218 528 219
rect 528 218 529 219
rect 529 218 530 219
rect 530 218 531 219
rect 531 218 532 219
rect 532 218 533 219
rect 90 217 91 218
rect 91 217 92 218
rect 92 217 93 218
rect 93 217 94 218
rect 94 217 95 218
rect 95 217 96 218
rect 96 217 97 218
rect 97 217 98 218
rect 98 217 99 218
rect 175 217 176 218
rect 176 217 177 218
rect 177 217 178 218
rect 178 217 179 218
rect 179 217 180 218
rect 180 217 181 218
rect 181 217 182 218
rect 182 217 183 218
rect 183 217 184 218
rect 184 217 185 218
rect 185 217 186 218
rect 186 217 187 218
rect 187 217 188 218
rect 188 217 189 218
rect 189 217 190 218
rect 190 217 191 218
rect 191 217 192 218
rect 192 217 193 218
rect 193 217 194 218
rect 194 217 195 218
rect 195 217 196 218
rect 196 217 197 218
rect 197 217 198 218
rect 198 217 199 218
rect 199 217 200 218
rect 200 217 201 218
rect 201 217 202 218
rect 202 217 203 218
rect 203 217 204 218
rect 204 217 205 218
rect 205 217 206 218
rect 206 217 207 218
rect 207 217 208 218
rect 208 217 209 218
rect 209 217 210 218
rect 210 217 211 218
rect 211 217 212 218
rect 212 217 213 218
rect 414 217 415 218
rect 415 217 416 218
rect 416 217 417 218
rect 435 217 436 218
rect 436 217 437 218
rect 437 217 438 218
rect 438 217 439 218
rect 439 217 440 218
rect 440 217 441 218
rect 441 217 442 218
rect 442 217 443 218
rect 443 217 444 218
rect 444 217 445 218
rect 461 217 462 218
rect 462 217 463 218
rect 463 217 464 218
rect 464 217 465 218
rect 465 217 466 218
rect 474 217 475 218
rect 475 217 476 218
rect 476 217 477 218
rect 477 217 478 218
rect 478 217 479 218
rect 479 217 480 218
rect 480 217 481 218
rect 481 217 482 218
rect 482 217 483 218
rect 483 217 484 218
rect 484 217 485 218
rect 485 217 486 218
rect 486 217 487 218
rect 487 217 488 218
rect 523 217 524 218
rect 524 217 525 218
rect 525 217 526 218
rect 526 217 527 218
rect 527 217 528 218
rect 528 217 529 218
rect 529 217 530 218
rect 530 217 531 218
rect 531 217 532 218
rect 532 217 533 218
rect 90 216 91 217
rect 91 216 92 217
rect 92 216 93 217
rect 93 216 94 217
rect 94 216 95 217
rect 95 216 96 217
rect 96 216 97 217
rect 97 216 98 217
rect 98 216 99 217
rect 175 216 176 217
rect 176 216 177 217
rect 177 216 178 217
rect 178 216 179 217
rect 179 216 180 217
rect 180 216 181 217
rect 181 216 182 217
rect 182 216 183 217
rect 183 216 184 217
rect 184 216 185 217
rect 185 216 186 217
rect 186 216 187 217
rect 187 216 188 217
rect 188 216 189 217
rect 189 216 190 217
rect 190 216 191 217
rect 191 216 192 217
rect 192 216 193 217
rect 193 216 194 217
rect 194 216 195 217
rect 195 216 196 217
rect 196 216 197 217
rect 197 216 198 217
rect 198 216 199 217
rect 199 216 200 217
rect 200 216 201 217
rect 201 216 202 217
rect 202 216 203 217
rect 203 216 204 217
rect 204 216 205 217
rect 205 216 206 217
rect 206 216 207 217
rect 207 216 208 217
rect 208 216 209 217
rect 209 216 210 217
rect 210 216 211 217
rect 211 216 212 217
rect 212 216 213 217
rect 414 216 415 217
rect 415 216 416 217
rect 416 216 417 217
rect 435 216 436 217
rect 436 216 437 217
rect 437 216 438 217
rect 438 216 439 217
rect 439 216 440 217
rect 440 216 441 217
rect 441 216 442 217
rect 442 216 443 217
rect 443 216 444 217
rect 444 216 445 217
rect 463 216 464 217
rect 464 216 465 217
rect 465 216 466 217
rect 474 216 475 217
rect 475 216 476 217
rect 476 216 477 217
rect 477 216 478 217
rect 478 216 479 217
rect 479 216 480 217
rect 480 216 481 217
rect 481 216 482 217
rect 482 216 483 217
rect 483 216 484 217
rect 484 216 485 217
rect 485 216 486 217
rect 486 216 487 217
rect 487 216 488 217
rect 523 216 524 217
rect 524 216 525 217
rect 525 216 526 217
rect 526 216 527 217
rect 527 216 528 217
rect 528 216 529 217
rect 529 216 530 217
rect 530 216 531 217
rect 531 216 532 217
rect 532 216 533 217
rect 90 215 91 216
rect 91 215 92 216
rect 92 215 93 216
rect 93 215 94 216
rect 94 215 95 216
rect 95 215 96 216
rect 96 215 97 216
rect 97 215 98 216
rect 98 215 99 216
rect 99 215 100 216
rect 100 215 101 216
rect 175 215 176 216
rect 176 215 177 216
rect 177 215 178 216
rect 178 215 179 216
rect 179 215 180 216
rect 180 215 181 216
rect 181 215 182 216
rect 182 215 183 216
rect 183 215 184 216
rect 184 215 185 216
rect 185 215 186 216
rect 186 215 187 216
rect 187 215 188 216
rect 188 215 189 216
rect 189 215 190 216
rect 190 215 191 216
rect 191 215 192 216
rect 192 215 193 216
rect 193 215 194 216
rect 194 215 195 216
rect 195 215 196 216
rect 196 215 197 216
rect 197 215 198 216
rect 198 215 199 216
rect 199 215 200 216
rect 200 215 201 216
rect 201 215 202 216
rect 202 215 203 216
rect 203 215 204 216
rect 204 215 205 216
rect 205 215 206 216
rect 206 215 207 216
rect 207 215 208 216
rect 208 215 209 216
rect 209 215 210 216
rect 210 215 211 216
rect 211 215 212 216
rect 212 215 213 216
rect 414 215 415 216
rect 415 215 416 216
rect 416 215 417 216
rect 435 215 436 216
rect 436 215 437 216
rect 437 215 438 216
rect 438 215 439 216
rect 439 215 440 216
rect 440 215 441 216
rect 441 215 442 216
rect 442 215 443 216
rect 443 215 444 216
rect 444 215 445 216
rect 463 215 464 216
rect 464 215 465 216
rect 465 215 466 216
rect 469 215 470 216
rect 470 215 471 216
rect 471 215 472 216
rect 472 215 473 216
rect 473 215 474 216
rect 474 215 475 216
rect 475 215 476 216
rect 476 215 477 216
rect 477 215 478 216
rect 478 215 479 216
rect 479 215 480 216
rect 480 215 481 216
rect 481 215 482 216
rect 482 215 483 216
rect 483 215 484 216
rect 484 215 485 216
rect 485 215 486 216
rect 486 215 487 216
rect 487 215 488 216
rect 488 215 489 216
rect 489 215 490 216
rect 490 215 491 216
rect 491 215 492 216
rect 492 215 493 216
rect 493 215 494 216
rect 494 215 495 216
rect 495 215 496 216
rect 523 215 524 216
rect 524 215 525 216
rect 525 215 526 216
rect 526 215 527 216
rect 527 215 528 216
rect 528 215 529 216
rect 529 215 530 216
rect 530 215 531 216
rect 531 215 532 216
rect 532 215 533 216
rect 90 214 91 215
rect 91 214 92 215
rect 92 214 93 215
rect 93 214 94 215
rect 94 214 95 215
rect 95 214 96 215
rect 96 214 97 215
rect 97 214 98 215
rect 98 214 99 215
rect 99 214 100 215
rect 100 214 101 215
rect 175 214 176 215
rect 176 214 177 215
rect 177 214 178 215
rect 178 214 179 215
rect 179 214 180 215
rect 180 214 181 215
rect 203 214 204 215
rect 204 214 205 215
rect 205 214 206 215
rect 206 214 207 215
rect 207 214 208 215
rect 208 214 209 215
rect 209 214 210 215
rect 210 214 211 215
rect 211 214 212 215
rect 212 214 213 215
rect 435 214 436 215
rect 436 214 437 215
rect 437 214 438 215
rect 438 214 439 215
rect 439 214 440 215
rect 440 214 441 215
rect 441 214 442 215
rect 442 214 443 215
rect 443 214 444 215
rect 444 214 445 215
rect 469 214 470 215
rect 470 214 471 215
rect 471 214 472 215
rect 472 214 473 215
rect 473 214 474 215
rect 474 214 475 215
rect 475 214 476 215
rect 476 214 477 215
rect 477 214 478 215
rect 478 214 479 215
rect 479 214 480 215
rect 480 214 481 215
rect 481 214 482 215
rect 482 214 483 215
rect 483 214 484 215
rect 484 214 485 215
rect 485 214 486 215
rect 486 214 487 215
rect 487 214 488 215
rect 488 214 489 215
rect 489 214 490 215
rect 490 214 491 215
rect 491 214 492 215
rect 492 214 493 215
rect 493 214 494 215
rect 494 214 495 215
rect 495 214 496 215
rect 523 214 524 215
rect 524 214 525 215
rect 525 214 526 215
rect 526 214 527 215
rect 527 214 528 215
rect 528 214 529 215
rect 529 214 530 215
rect 530 214 531 215
rect 531 214 532 215
rect 532 214 533 215
rect 90 213 91 214
rect 91 213 92 214
rect 92 213 93 214
rect 93 213 94 214
rect 94 213 95 214
rect 95 213 96 214
rect 96 213 97 214
rect 97 213 98 214
rect 98 213 99 214
rect 99 213 100 214
rect 100 213 101 214
rect 173 213 174 214
rect 174 213 175 214
rect 175 213 176 214
rect 176 213 177 214
rect 177 213 178 214
rect 178 213 179 214
rect 179 213 180 214
rect 180 213 181 214
rect 203 213 204 214
rect 204 213 205 214
rect 205 213 206 214
rect 206 213 207 214
rect 207 213 208 214
rect 208 213 209 214
rect 209 213 210 214
rect 210 213 211 214
rect 211 213 212 214
rect 212 213 213 214
rect 213 213 214 214
rect 214 213 215 214
rect 433 213 434 214
rect 434 213 435 214
rect 435 213 436 214
rect 436 213 437 214
rect 437 213 438 214
rect 438 213 439 214
rect 439 213 440 214
rect 440 213 441 214
rect 441 213 442 214
rect 442 213 443 214
rect 443 213 444 214
rect 444 213 445 214
rect 469 213 470 214
rect 470 213 471 214
rect 471 213 472 214
rect 472 213 473 214
rect 473 213 474 214
rect 474 213 475 214
rect 475 213 476 214
rect 476 213 477 214
rect 477 213 478 214
rect 478 213 479 214
rect 479 213 480 214
rect 480 213 481 214
rect 481 213 482 214
rect 482 213 483 214
rect 483 213 484 214
rect 484 213 485 214
rect 485 213 486 214
rect 486 213 487 214
rect 487 213 488 214
rect 488 213 489 214
rect 489 213 490 214
rect 490 213 491 214
rect 491 213 492 214
rect 492 213 493 214
rect 493 213 494 214
rect 494 213 495 214
rect 495 213 496 214
rect 521 213 522 214
rect 522 213 523 214
rect 523 213 524 214
rect 524 213 525 214
rect 525 213 526 214
rect 526 213 527 214
rect 527 213 528 214
rect 528 213 529 214
rect 529 213 530 214
rect 530 213 531 214
rect 531 213 532 214
rect 532 213 533 214
rect 90 212 91 213
rect 91 212 92 213
rect 92 212 93 213
rect 93 212 94 213
rect 94 212 95 213
rect 95 212 96 213
rect 96 212 97 213
rect 97 212 98 213
rect 98 212 99 213
rect 99 212 100 213
rect 100 212 101 213
rect 173 212 174 213
rect 174 212 175 213
rect 175 212 176 213
rect 176 212 177 213
rect 177 212 178 213
rect 178 212 179 213
rect 203 212 204 213
rect 204 212 205 213
rect 205 212 206 213
rect 206 212 207 213
rect 207 212 208 213
rect 208 212 209 213
rect 209 212 210 213
rect 210 212 211 213
rect 211 212 212 213
rect 212 212 213 213
rect 213 212 214 213
rect 214 212 215 213
rect 433 212 434 213
rect 434 212 435 213
rect 435 212 436 213
rect 436 212 437 213
rect 437 212 438 213
rect 438 212 439 213
rect 439 212 440 213
rect 440 212 441 213
rect 441 212 442 213
rect 442 212 443 213
rect 443 212 444 213
rect 444 212 445 213
rect 469 212 470 213
rect 470 212 471 213
rect 471 212 472 213
rect 474 212 475 213
rect 475 212 476 213
rect 476 212 477 213
rect 480 212 481 213
rect 481 212 482 213
rect 482 212 483 213
rect 487 212 488 213
rect 488 212 489 213
rect 489 212 490 213
rect 491 212 492 213
rect 492 212 493 213
rect 493 212 494 213
rect 521 212 522 213
rect 522 212 523 213
rect 523 212 524 213
rect 524 212 525 213
rect 525 212 526 213
rect 526 212 527 213
rect 527 212 528 213
rect 528 212 529 213
rect 529 212 530 213
rect 530 212 531 213
rect 531 212 532 213
rect 532 212 533 213
rect 90 211 91 212
rect 91 211 92 212
rect 92 211 93 212
rect 93 211 94 212
rect 94 211 95 212
rect 95 211 96 212
rect 96 211 97 212
rect 97 211 98 212
rect 98 211 99 212
rect 99 211 100 212
rect 100 211 101 212
rect 173 211 174 212
rect 174 211 175 212
rect 175 211 176 212
rect 176 211 177 212
rect 177 211 178 212
rect 178 211 179 212
rect 203 211 204 212
rect 204 211 205 212
rect 205 211 206 212
rect 206 211 207 212
rect 207 211 208 212
rect 208 211 209 212
rect 209 211 210 212
rect 210 211 211 212
rect 211 211 212 212
rect 212 211 213 212
rect 213 211 214 212
rect 214 211 215 212
rect 433 211 434 212
rect 434 211 435 212
rect 435 211 436 212
rect 436 211 437 212
rect 437 211 438 212
rect 438 211 439 212
rect 439 211 440 212
rect 440 211 441 212
rect 441 211 442 212
rect 442 211 443 212
rect 443 211 444 212
rect 444 211 445 212
rect 469 211 470 212
rect 470 211 471 212
rect 471 211 472 212
rect 474 211 475 212
rect 475 211 476 212
rect 476 211 477 212
rect 480 211 481 212
rect 481 211 482 212
rect 482 211 483 212
rect 487 211 488 212
rect 488 211 489 212
rect 489 211 490 212
rect 491 211 492 212
rect 492 211 493 212
rect 493 211 494 212
rect 521 211 522 212
rect 522 211 523 212
rect 523 211 524 212
rect 524 211 525 212
rect 525 211 526 212
rect 526 211 527 212
rect 527 211 528 212
rect 528 211 529 212
rect 529 211 530 212
rect 530 211 531 212
rect 531 211 532 212
rect 532 211 533 212
rect 92 210 93 211
rect 93 210 94 211
rect 94 210 95 211
rect 95 210 96 211
rect 96 210 97 211
rect 97 210 98 211
rect 98 210 99 211
rect 99 210 100 211
rect 100 210 101 211
rect 173 210 174 211
rect 174 210 175 211
rect 175 210 176 211
rect 176 210 177 211
rect 177 210 178 211
rect 178 210 179 211
rect 205 210 206 211
rect 206 210 207 211
rect 207 210 208 211
rect 208 210 209 211
rect 209 210 210 211
rect 210 210 211 211
rect 211 210 212 211
rect 212 210 213 211
rect 213 210 214 211
rect 214 210 215 211
rect 435 210 436 211
rect 436 210 437 211
rect 437 210 438 211
rect 438 210 439 211
rect 439 210 440 211
rect 440 210 441 211
rect 441 210 442 211
rect 442 210 443 211
rect 443 210 444 211
rect 444 210 445 211
rect 521 210 522 211
rect 522 210 523 211
rect 523 210 524 211
rect 524 210 525 211
rect 525 210 526 211
rect 526 210 527 211
rect 527 210 528 211
rect 528 210 529 211
rect 529 210 530 211
rect 530 210 531 211
rect 92 209 93 210
rect 93 209 94 210
rect 94 209 95 210
rect 95 209 96 210
rect 96 209 97 210
rect 97 209 98 210
rect 98 209 99 210
rect 99 209 100 210
rect 100 209 101 210
rect 101 209 102 210
rect 102 209 103 210
rect 173 209 174 210
rect 174 209 175 210
rect 175 209 176 210
rect 176 209 177 210
rect 177 209 178 210
rect 178 209 179 210
rect 205 209 206 210
rect 206 209 207 210
rect 207 209 208 210
rect 208 209 209 210
rect 209 209 210 210
rect 210 209 211 210
rect 211 209 212 210
rect 212 209 213 210
rect 213 209 214 210
rect 214 209 215 210
rect 215 209 216 210
rect 216 209 217 210
rect 435 209 436 210
rect 436 209 437 210
rect 437 209 438 210
rect 438 209 439 210
rect 439 209 440 210
rect 440 209 441 210
rect 441 209 442 210
rect 442 209 443 210
rect 443 209 444 210
rect 444 209 445 210
rect 521 209 522 210
rect 522 209 523 210
rect 523 209 524 210
rect 524 209 525 210
rect 525 209 526 210
rect 526 209 527 210
rect 527 209 528 210
rect 528 209 529 210
rect 529 209 530 210
rect 530 209 531 210
rect 92 208 93 209
rect 93 208 94 209
rect 94 208 95 209
rect 95 208 96 209
rect 96 208 97 209
rect 97 208 98 209
rect 98 208 99 209
rect 99 208 100 209
rect 100 208 101 209
rect 101 208 102 209
rect 102 208 103 209
rect 173 208 174 209
rect 174 208 175 209
rect 175 208 176 209
rect 176 208 177 209
rect 177 208 178 209
rect 178 208 179 209
rect 205 208 206 209
rect 206 208 207 209
rect 207 208 208 209
rect 208 208 209 209
rect 209 208 210 209
rect 210 208 211 209
rect 211 208 212 209
rect 212 208 213 209
rect 213 208 214 209
rect 214 208 215 209
rect 215 208 216 209
rect 216 208 217 209
rect 435 208 436 209
rect 436 208 437 209
rect 437 208 438 209
rect 438 208 439 209
rect 439 208 440 209
rect 440 208 441 209
rect 441 208 442 209
rect 442 208 443 209
rect 443 208 444 209
rect 444 208 445 209
rect 521 208 522 209
rect 522 208 523 209
rect 523 208 524 209
rect 524 208 525 209
rect 525 208 526 209
rect 526 208 527 209
rect 527 208 528 209
rect 528 208 529 209
rect 529 208 530 209
rect 530 208 531 209
rect 92 207 93 208
rect 93 207 94 208
rect 94 207 95 208
rect 95 207 96 208
rect 96 207 97 208
rect 97 207 98 208
rect 98 207 99 208
rect 99 207 100 208
rect 100 207 101 208
rect 101 207 102 208
rect 102 207 103 208
rect 171 207 172 208
rect 172 207 173 208
rect 173 207 174 208
rect 174 207 175 208
rect 175 207 176 208
rect 176 207 177 208
rect 177 207 178 208
rect 178 207 179 208
rect 205 207 206 208
rect 206 207 207 208
rect 207 207 208 208
rect 208 207 209 208
rect 209 207 210 208
rect 210 207 211 208
rect 211 207 212 208
rect 212 207 213 208
rect 213 207 214 208
rect 214 207 215 208
rect 215 207 216 208
rect 216 207 217 208
rect 433 207 434 208
rect 434 207 435 208
rect 435 207 436 208
rect 436 207 437 208
rect 437 207 438 208
rect 438 207 439 208
rect 439 207 440 208
rect 440 207 441 208
rect 441 207 442 208
rect 442 207 443 208
rect 443 207 444 208
rect 444 207 445 208
rect 519 207 520 208
rect 520 207 521 208
rect 521 207 522 208
rect 522 207 523 208
rect 523 207 524 208
rect 524 207 525 208
rect 525 207 526 208
rect 526 207 527 208
rect 527 207 528 208
rect 528 207 529 208
rect 529 207 530 208
rect 530 207 531 208
rect 92 206 93 207
rect 93 206 94 207
rect 94 206 95 207
rect 95 206 96 207
rect 96 206 97 207
rect 97 206 98 207
rect 98 206 99 207
rect 99 206 100 207
rect 100 206 101 207
rect 101 206 102 207
rect 102 206 103 207
rect 171 206 172 207
rect 172 206 173 207
rect 173 206 174 207
rect 174 206 175 207
rect 175 206 176 207
rect 176 206 177 207
rect 206 206 207 207
rect 207 206 208 207
rect 208 206 209 207
rect 209 206 210 207
rect 210 206 211 207
rect 211 206 212 207
rect 212 206 213 207
rect 213 206 214 207
rect 214 206 215 207
rect 215 206 216 207
rect 216 206 217 207
rect 433 206 434 207
rect 434 206 435 207
rect 435 206 436 207
rect 436 206 437 207
rect 437 206 438 207
rect 438 206 439 207
rect 439 206 440 207
rect 440 206 441 207
rect 441 206 442 207
rect 442 206 443 207
rect 443 206 444 207
rect 444 206 445 207
rect 519 206 520 207
rect 520 206 521 207
rect 521 206 522 207
rect 522 206 523 207
rect 523 206 524 207
rect 524 206 525 207
rect 525 206 526 207
rect 526 206 527 207
rect 527 206 528 207
rect 528 206 529 207
rect 529 206 530 207
rect 530 206 531 207
rect 92 205 93 206
rect 93 205 94 206
rect 94 205 95 206
rect 95 205 96 206
rect 96 205 97 206
rect 97 205 98 206
rect 98 205 99 206
rect 99 205 100 206
rect 100 205 101 206
rect 101 205 102 206
rect 102 205 103 206
rect 171 205 172 206
rect 172 205 173 206
rect 173 205 174 206
rect 174 205 175 206
rect 175 205 176 206
rect 176 205 177 206
rect 206 205 207 206
rect 207 205 208 206
rect 208 205 209 206
rect 209 205 210 206
rect 210 205 211 206
rect 211 205 212 206
rect 212 205 213 206
rect 213 205 214 206
rect 214 205 215 206
rect 215 205 216 206
rect 216 205 217 206
rect 217 205 218 206
rect 218 205 219 206
rect 225 205 226 206
rect 226 205 227 206
rect 227 205 228 206
rect 228 205 229 206
rect 229 205 230 206
rect 433 205 434 206
rect 434 205 435 206
rect 435 205 436 206
rect 436 205 437 206
rect 437 205 438 206
rect 438 205 439 206
rect 439 205 440 206
rect 440 205 441 206
rect 441 205 442 206
rect 442 205 443 206
rect 443 205 444 206
rect 444 205 445 206
rect 519 205 520 206
rect 520 205 521 206
rect 521 205 522 206
rect 522 205 523 206
rect 523 205 524 206
rect 524 205 525 206
rect 525 205 526 206
rect 526 205 527 206
rect 527 205 528 206
rect 528 205 529 206
rect 529 205 530 206
rect 530 205 531 206
rect 92 204 93 205
rect 93 204 94 205
rect 94 204 95 205
rect 95 204 96 205
rect 96 204 97 205
rect 97 204 98 205
rect 98 204 99 205
rect 99 204 100 205
rect 100 204 101 205
rect 101 204 102 205
rect 102 204 103 205
rect 171 204 172 205
rect 172 204 173 205
rect 173 204 174 205
rect 174 204 175 205
rect 175 204 176 205
rect 176 204 177 205
rect 206 204 207 205
rect 207 204 208 205
rect 208 204 209 205
rect 209 204 210 205
rect 210 204 211 205
rect 211 204 212 205
rect 212 204 213 205
rect 213 204 214 205
rect 214 204 215 205
rect 215 204 216 205
rect 216 204 217 205
rect 217 204 218 205
rect 218 204 219 205
rect 225 204 226 205
rect 226 204 227 205
rect 227 204 228 205
rect 228 204 229 205
rect 229 204 230 205
rect 435 204 436 205
rect 436 204 437 205
rect 437 204 438 205
rect 438 204 439 205
rect 439 204 440 205
rect 440 204 441 205
rect 441 204 442 205
rect 442 204 443 205
rect 443 204 444 205
rect 444 204 445 205
rect 519 204 520 205
rect 520 204 521 205
rect 521 204 522 205
rect 522 204 523 205
rect 523 204 524 205
rect 524 204 525 205
rect 525 204 526 205
rect 526 204 527 205
rect 527 204 528 205
rect 528 204 529 205
rect 529 204 530 205
rect 92 203 93 204
rect 93 203 94 204
rect 94 203 95 204
rect 95 203 96 204
rect 96 203 97 204
rect 97 203 98 204
rect 98 203 99 204
rect 99 203 100 204
rect 100 203 101 204
rect 101 203 102 204
rect 102 203 103 204
rect 169 203 170 204
rect 170 203 171 204
rect 171 203 172 204
rect 172 203 173 204
rect 173 203 174 204
rect 174 203 175 204
rect 175 203 176 204
rect 176 203 177 204
rect 206 203 207 204
rect 207 203 208 204
rect 208 203 209 204
rect 209 203 210 204
rect 210 203 211 204
rect 211 203 212 204
rect 212 203 213 204
rect 213 203 214 204
rect 214 203 215 204
rect 215 203 216 204
rect 216 203 217 204
rect 217 203 218 204
rect 218 203 219 204
rect 225 203 226 204
rect 226 203 227 204
rect 227 203 228 204
rect 228 203 229 204
rect 229 203 230 204
rect 435 203 436 204
rect 436 203 437 204
rect 437 203 438 204
rect 438 203 439 204
rect 439 203 440 204
rect 440 203 441 204
rect 441 203 442 204
rect 442 203 443 204
rect 443 203 444 204
rect 444 203 445 204
rect 517 203 518 204
rect 518 203 519 204
rect 519 203 520 204
rect 520 203 521 204
rect 521 203 522 204
rect 522 203 523 204
rect 523 203 524 204
rect 524 203 525 204
rect 525 203 526 204
rect 526 203 527 204
rect 527 203 528 204
rect 528 203 529 204
rect 529 203 530 204
rect 94 202 95 203
rect 95 202 96 203
rect 96 202 97 203
rect 97 202 98 203
rect 98 202 99 203
rect 99 202 100 203
rect 100 202 101 203
rect 101 202 102 203
rect 102 202 103 203
rect 169 202 170 203
rect 170 202 171 203
rect 171 202 172 203
rect 172 202 173 203
rect 173 202 174 203
rect 174 202 175 203
rect 175 202 176 203
rect 206 202 207 203
rect 207 202 208 203
rect 208 202 209 203
rect 209 202 210 203
rect 210 202 211 203
rect 211 202 212 203
rect 212 202 213 203
rect 213 202 214 203
rect 214 202 215 203
rect 215 202 216 203
rect 216 202 217 203
rect 217 202 218 203
rect 218 202 219 203
rect 225 202 226 203
rect 226 202 227 203
rect 227 202 228 203
rect 228 202 229 203
rect 229 202 230 203
rect 435 202 436 203
rect 436 202 437 203
rect 437 202 438 203
rect 438 202 439 203
rect 439 202 440 203
rect 440 202 441 203
rect 441 202 442 203
rect 442 202 443 203
rect 443 202 444 203
rect 444 202 445 203
rect 517 202 518 203
rect 518 202 519 203
rect 519 202 520 203
rect 520 202 521 203
rect 521 202 522 203
rect 522 202 523 203
rect 523 202 524 203
rect 524 202 525 203
rect 525 202 526 203
rect 526 202 527 203
rect 527 202 528 203
rect 528 202 529 203
rect 529 202 530 203
rect 94 201 95 202
rect 95 201 96 202
rect 96 201 97 202
rect 97 201 98 202
rect 98 201 99 202
rect 99 201 100 202
rect 100 201 101 202
rect 101 201 102 202
rect 102 201 103 202
rect 169 201 170 202
rect 170 201 171 202
rect 171 201 172 202
rect 172 201 173 202
rect 173 201 174 202
rect 174 201 175 202
rect 175 201 176 202
rect 206 201 207 202
rect 207 201 208 202
rect 208 201 209 202
rect 209 201 210 202
rect 210 201 211 202
rect 211 201 212 202
rect 212 201 213 202
rect 213 201 214 202
rect 214 201 215 202
rect 215 201 216 202
rect 216 201 217 202
rect 217 201 218 202
rect 218 201 219 202
rect 225 201 226 202
rect 226 201 227 202
rect 227 201 228 202
rect 228 201 229 202
rect 229 201 230 202
rect 433 201 434 202
rect 434 201 435 202
rect 435 201 436 202
rect 436 201 437 202
rect 437 201 438 202
rect 438 201 439 202
rect 439 201 440 202
rect 440 201 441 202
rect 441 201 442 202
rect 442 201 443 202
rect 443 201 444 202
rect 444 201 445 202
rect 517 201 518 202
rect 518 201 519 202
rect 519 201 520 202
rect 520 201 521 202
rect 521 201 522 202
rect 522 201 523 202
rect 523 201 524 202
rect 524 201 525 202
rect 525 201 526 202
rect 526 201 527 202
rect 527 201 528 202
rect 528 201 529 202
rect 529 201 530 202
rect 94 200 95 201
rect 95 200 96 201
rect 96 200 97 201
rect 97 200 98 201
rect 98 200 99 201
rect 99 200 100 201
rect 100 200 101 201
rect 101 200 102 201
rect 102 200 103 201
rect 169 200 170 201
rect 170 200 171 201
rect 171 200 172 201
rect 172 200 173 201
rect 173 200 174 201
rect 174 200 175 201
rect 175 200 176 201
rect 206 200 207 201
rect 207 200 208 201
rect 208 200 209 201
rect 209 200 210 201
rect 210 200 211 201
rect 211 200 212 201
rect 212 200 213 201
rect 213 200 214 201
rect 214 200 215 201
rect 215 200 216 201
rect 216 200 217 201
rect 217 200 218 201
rect 218 200 219 201
rect 225 200 226 201
rect 226 200 227 201
rect 227 200 228 201
rect 228 200 229 201
rect 229 200 230 201
rect 433 200 434 201
rect 434 200 435 201
rect 435 200 436 201
rect 436 200 437 201
rect 437 200 438 201
rect 438 200 439 201
rect 439 200 440 201
rect 440 200 441 201
rect 441 200 442 201
rect 442 200 443 201
rect 443 200 444 201
rect 444 200 445 201
rect 517 200 518 201
rect 518 200 519 201
rect 519 200 520 201
rect 520 200 521 201
rect 521 200 522 201
rect 522 200 523 201
rect 523 200 524 201
rect 524 200 525 201
rect 525 200 526 201
rect 526 200 527 201
rect 527 200 528 201
rect 528 200 529 201
rect 529 200 530 201
rect 94 199 95 200
rect 95 199 96 200
rect 96 199 97 200
rect 97 199 98 200
rect 98 199 99 200
rect 99 199 100 200
rect 100 199 101 200
rect 101 199 102 200
rect 102 199 103 200
rect 103 199 104 200
rect 167 199 168 200
rect 168 199 169 200
rect 169 199 170 200
rect 170 199 171 200
rect 171 199 172 200
rect 172 199 173 200
rect 173 199 174 200
rect 174 199 175 200
rect 175 199 176 200
rect 176 199 177 200
rect 206 199 207 200
rect 207 199 208 200
rect 208 199 209 200
rect 209 199 210 200
rect 210 199 211 200
rect 211 199 212 200
rect 212 199 213 200
rect 213 199 214 200
rect 214 199 215 200
rect 215 199 216 200
rect 216 199 217 200
rect 217 199 218 200
rect 218 199 219 200
rect 219 199 220 200
rect 220 199 221 200
rect 223 199 224 200
rect 224 199 225 200
rect 225 199 226 200
rect 226 199 227 200
rect 227 199 228 200
rect 228 199 229 200
rect 229 199 230 200
rect 230 199 231 200
rect 231 199 232 200
rect 433 199 434 200
rect 434 199 435 200
rect 435 199 436 200
rect 436 199 437 200
rect 437 199 438 200
rect 438 199 439 200
rect 439 199 440 200
rect 440 199 441 200
rect 441 199 442 200
rect 442 199 443 200
rect 443 199 444 200
rect 444 199 445 200
rect 515 199 516 200
rect 516 199 517 200
rect 517 199 518 200
rect 518 199 519 200
rect 519 199 520 200
rect 520 199 521 200
rect 521 199 522 200
rect 522 199 523 200
rect 523 199 524 200
rect 524 199 525 200
rect 525 199 526 200
rect 526 199 527 200
rect 527 199 528 200
rect 528 199 529 200
rect 529 199 530 200
rect 94 198 95 199
rect 95 198 96 199
rect 96 198 97 199
rect 97 198 98 199
rect 98 198 99 199
rect 99 198 100 199
rect 100 198 101 199
rect 101 198 102 199
rect 102 198 103 199
rect 103 198 104 199
rect 167 198 168 199
rect 168 198 169 199
rect 169 198 170 199
rect 170 198 171 199
rect 171 198 172 199
rect 172 198 173 199
rect 173 198 174 199
rect 174 198 175 199
rect 175 198 176 199
rect 176 198 177 199
rect 206 198 207 199
rect 207 198 208 199
rect 208 198 209 199
rect 209 198 210 199
rect 210 198 211 199
rect 211 198 212 199
rect 212 198 213 199
rect 213 198 214 199
rect 214 198 215 199
rect 215 198 216 199
rect 216 198 217 199
rect 217 198 218 199
rect 218 198 219 199
rect 219 198 220 199
rect 220 198 221 199
rect 223 198 224 199
rect 224 198 225 199
rect 225 198 226 199
rect 226 198 227 199
rect 227 198 228 199
rect 228 198 229 199
rect 229 198 230 199
rect 230 198 231 199
rect 231 198 232 199
rect 435 198 436 199
rect 436 198 437 199
rect 437 198 438 199
rect 438 198 439 199
rect 439 198 440 199
rect 440 198 441 199
rect 441 198 442 199
rect 442 198 443 199
rect 443 198 444 199
rect 444 198 445 199
rect 515 198 516 199
rect 516 198 517 199
rect 517 198 518 199
rect 518 198 519 199
rect 519 198 520 199
rect 520 198 521 199
rect 521 198 522 199
rect 522 198 523 199
rect 523 198 524 199
rect 524 198 525 199
rect 525 198 526 199
rect 526 198 527 199
rect 527 198 528 199
rect 528 198 529 199
rect 529 198 530 199
rect 94 197 95 198
rect 95 197 96 198
rect 96 197 97 198
rect 97 197 98 198
rect 98 197 99 198
rect 99 197 100 198
rect 100 197 101 198
rect 101 197 102 198
rect 102 197 103 198
rect 103 197 104 198
rect 163 197 164 198
rect 164 197 165 198
rect 165 197 166 198
rect 166 197 167 198
rect 167 197 168 198
rect 168 197 169 198
rect 169 197 170 198
rect 170 197 171 198
rect 171 197 172 198
rect 172 197 173 198
rect 173 197 174 198
rect 174 197 175 198
rect 175 197 176 198
rect 176 197 177 198
rect 177 197 178 198
rect 178 197 179 198
rect 179 197 180 198
rect 180 197 181 198
rect 201 197 202 198
rect 202 197 203 198
rect 203 197 204 198
rect 205 197 206 198
rect 206 197 207 198
rect 207 197 208 198
rect 208 197 209 198
rect 209 197 210 198
rect 210 197 211 198
rect 211 197 212 198
rect 212 197 213 198
rect 213 197 214 198
rect 214 197 215 198
rect 215 197 216 198
rect 216 197 217 198
rect 217 197 218 198
rect 218 197 219 198
rect 219 197 220 198
rect 220 197 221 198
rect 221 197 222 198
rect 223 197 224 198
rect 224 197 225 198
rect 225 197 226 198
rect 226 197 227 198
rect 227 197 228 198
rect 228 197 229 198
rect 229 197 230 198
rect 230 197 231 198
rect 231 197 232 198
rect 360 197 361 198
rect 361 197 362 198
rect 362 197 363 198
rect 363 197 364 198
rect 364 197 365 198
rect 365 197 366 198
rect 366 197 367 198
rect 367 197 368 198
rect 368 197 369 198
rect 369 197 370 198
rect 370 197 371 198
rect 371 197 372 198
rect 372 197 373 198
rect 373 197 374 198
rect 374 197 375 198
rect 375 197 376 198
rect 376 197 377 198
rect 377 197 378 198
rect 378 197 379 198
rect 379 197 380 198
rect 380 197 381 198
rect 381 197 382 198
rect 382 197 383 198
rect 383 197 384 198
rect 384 197 385 198
rect 385 197 386 198
rect 386 197 387 198
rect 387 197 388 198
rect 388 197 389 198
rect 390 197 391 198
rect 391 197 392 198
rect 392 197 393 198
rect 393 197 394 198
rect 394 197 395 198
rect 395 197 396 198
rect 396 197 397 198
rect 397 197 398 198
rect 398 197 399 198
rect 399 197 400 198
rect 400 197 401 198
rect 401 197 402 198
rect 402 197 403 198
rect 403 197 404 198
rect 404 197 405 198
rect 405 197 406 198
rect 406 197 407 198
rect 407 197 408 198
rect 435 197 436 198
rect 436 197 437 198
rect 437 197 438 198
rect 438 197 439 198
rect 439 197 440 198
rect 440 197 441 198
rect 441 197 442 198
rect 442 197 443 198
rect 443 197 444 198
rect 444 197 445 198
rect 515 197 516 198
rect 516 197 517 198
rect 517 197 518 198
rect 518 197 519 198
rect 519 197 520 198
rect 520 197 521 198
rect 521 197 522 198
rect 522 197 523 198
rect 523 197 524 198
rect 524 197 525 198
rect 525 197 526 198
rect 526 197 527 198
rect 527 197 528 198
rect 528 197 529 198
rect 529 197 530 198
rect 94 196 95 197
rect 95 196 96 197
rect 96 196 97 197
rect 97 196 98 197
rect 98 196 99 197
rect 99 196 100 197
rect 100 196 101 197
rect 101 196 102 197
rect 102 196 103 197
rect 103 196 104 197
rect 163 196 164 197
rect 164 196 165 197
rect 165 196 166 197
rect 166 196 167 197
rect 167 196 168 197
rect 168 196 169 197
rect 169 196 170 197
rect 170 196 171 197
rect 171 196 172 197
rect 172 196 173 197
rect 173 196 174 197
rect 174 196 175 197
rect 175 196 176 197
rect 176 196 177 197
rect 177 196 178 197
rect 178 196 179 197
rect 179 196 180 197
rect 180 196 181 197
rect 201 196 202 197
rect 202 196 203 197
rect 203 196 204 197
rect 205 196 206 197
rect 206 196 207 197
rect 207 196 208 197
rect 208 196 209 197
rect 209 196 210 197
rect 210 196 211 197
rect 211 196 212 197
rect 212 196 213 197
rect 213 196 214 197
rect 214 196 215 197
rect 215 196 216 197
rect 216 196 217 197
rect 217 196 218 197
rect 218 196 219 197
rect 219 196 220 197
rect 220 196 221 197
rect 221 196 222 197
rect 223 196 224 197
rect 224 196 225 197
rect 225 196 226 197
rect 226 196 227 197
rect 227 196 228 197
rect 228 196 229 197
rect 229 196 230 197
rect 230 196 231 197
rect 231 196 232 197
rect 360 196 361 197
rect 361 196 362 197
rect 362 196 363 197
rect 363 196 364 197
rect 364 196 365 197
rect 365 196 366 197
rect 366 196 367 197
rect 367 196 368 197
rect 368 196 369 197
rect 369 196 370 197
rect 370 196 371 197
rect 371 196 372 197
rect 372 196 373 197
rect 373 196 374 197
rect 374 196 375 197
rect 375 196 376 197
rect 376 196 377 197
rect 377 196 378 197
rect 378 196 379 197
rect 379 196 380 197
rect 380 196 381 197
rect 381 196 382 197
rect 382 196 383 197
rect 383 196 384 197
rect 384 196 385 197
rect 385 196 386 197
rect 386 196 387 197
rect 387 196 388 197
rect 388 196 389 197
rect 390 196 391 197
rect 391 196 392 197
rect 392 196 393 197
rect 393 196 394 197
rect 394 196 395 197
rect 395 196 396 197
rect 396 196 397 197
rect 397 196 398 197
rect 398 196 399 197
rect 399 196 400 197
rect 400 196 401 197
rect 401 196 402 197
rect 402 196 403 197
rect 403 196 404 197
rect 404 196 405 197
rect 405 196 406 197
rect 406 196 407 197
rect 407 196 408 197
rect 435 196 436 197
rect 436 196 437 197
rect 437 196 438 197
rect 438 196 439 197
rect 439 196 440 197
rect 440 196 441 197
rect 441 196 442 197
rect 442 196 443 197
rect 443 196 444 197
rect 444 196 445 197
rect 515 196 516 197
rect 516 196 517 197
rect 517 196 518 197
rect 518 196 519 197
rect 519 196 520 197
rect 520 196 521 197
rect 521 196 522 197
rect 522 196 523 197
rect 523 196 524 197
rect 524 196 525 197
rect 525 196 526 197
rect 526 196 527 197
rect 527 196 528 197
rect 94 195 95 196
rect 95 195 96 196
rect 96 195 97 196
rect 97 195 98 196
rect 98 195 99 196
rect 99 195 100 196
rect 100 195 101 196
rect 101 195 102 196
rect 102 195 103 196
rect 103 195 104 196
rect 163 195 164 196
rect 164 195 165 196
rect 165 195 166 196
rect 166 195 167 196
rect 167 195 168 196
rect 168 195 169 196
rect 169 195 170 196
rect 170 195 171 196
rect 171 195 172 196
rect 172 195 173 196
rect 173 195 174 196
rect 174 195 175 196
rect 175 195 176 196
rect 176 195 177 196
rect 177 195 178 196
rect 178 195 179 196
rect 179 195 180 196
rect 180 195 181 196
rect 201 195 202 196
rect 202 195 203 196
rect 203 195 204 196
rect 204 195 205 196
rect 205 195 206 196
rect 206 195 207 196
rect 207 195 208 196
rect 208 195 209 196
rect 209 195 210 196
rect 210 195 211 196
rect 211 195 212 196
rect 212 195 213 196
rect 213 195 214 196
rect 214 195 215 196
rect 215 195 216 196
rect 216 195 217 196
rect 217 195 218 196
rect 218 195 219 196
rect 219 195 220 196
rect 220 195 221 196
rect 221 195 222 196
rect 222 195 223 196
rect 223 195 224 196
rect 224 195 225 196
rect 225 195 226 196
rect 226 195 227 196
rect 227 195 228 196
rect 228 195 229 196
rect 229 195 230 196
rect 230 195 231 196
rect 231 195 232 196
rect 232 195 233 196
rect 233 195 234 196
rect 360 195 361 196
rect 361 195 362 196
rect 362 195 363 196
rect 363 195 364 196
rect 364 195 365 196
rect 365 195 366 196
rect 366 195 367 196
rect 367 195 368 196
rect 368 195 369 196
rect 369 195 370 196
rect 370 195 371 196
rect 371 195 372 196
rect 372 195 373 196
rect 373 195 374 196
rect 374 195 375 196
rect 375 195 376 196
rect 376 195 377 196
rect 377 195 378 196
rect 378 195 379 196
rect 379 195 380 196
rect 380 195 381 196
rect 381 195 382 196
rect 382 195 383 196
rect 383 195 384 196
rect 384 195 385 196
rect 385 195 386 196
rect 386 195 387 196
rect 387 195 388 196
rect 388 195 389 196
rect 389 195 390 196
rect 390 195 391 196
rect 391 195 392 196
rect 392 195 393 196
rect 393 195 394 196
rect 394 195 395 196
rect 395 195 396 196
rect 396 195 397 196
rect 397 195 398 196
rect 398 195 399 196
rect 399 195 400 196
rect 400 195 401 196
rect 401 195 402 196
rect 402 195 403 196
rect 403 195 404 196
rect 404 195 405 196
rect 405 195 406 196
rect 406 195 407 196
rect 407 195 408 196
rect 433 195 434 196
rect 434 195 435 196
rect 435 195 436 196
rect 436 195 437 196
rect 437 195 438 196
rect 438 195 439 196
rect 439 195 440 196
rect 440 195 441 196
rect 441 195 442 196
rect 442 195 443 196
rect 443 195 444 196
rect 444 195 445 196
rect 514 195 515 196
rect 515 195 516 196
rect 516 195 517 196
rect 517 195 518 196
rect 518 195 519 196
rect 519 195 520 196
rect 520 195 521 196
rect 521 195 522 196
rect 522 195 523 196
rect 523 195 524 196
rect 524 195 525 196
rect 525 195 526 196
rect 526 195 527 196
rect 527 195 528 196
rect 94 194 95 195
rect 95 194 96 195
rect 96 194 97 195
rect 97 194 98 195
rect 98 194 99 195
rect 99 194 100 195
rect 100 194 101 195
rect 101 194 102 195
rect 102 194 103 195
rect 103 194 104 195
rect 165 194 166 195
rect 166 194 167 195
rect 167 194 168 195
rect 169 194 170 195
rect 170 194 171 195
rect 171 194 172 195
rect 172 194 173 195
rect 173 194 174 195
rect 174 194 175 195
rect 175 194 176 195
rect 176 194 177 195
rect 177 194 178 195
rect 178 194 179 195
rect 179 194 180 195
rect 180 194 181 195
rect 203 194 204 195
rect 204 194 205 195
rect 205 194 206 195
rect 206 194 207 195
rect 208 194 209 195
rect 209 194 210 195
rect 210 194 211 195
rect 211 194 212 195
rect 212 194 213 195
rect 214 194 215 195
rect 215 194 216 195
rect 216 194 217 195
rect 217 194 218 195
rect 218 194 219 195
rect 220 194 221 195
rect 221 194 222 195
rect 222 194 223 195
rect 223 194 224 195
rect 224 194 225 195
rect 225 194 226 195
rect 226 194 227 195
rect 227 194 228 195
rect 228 194 229 195
rect 229 194 230 195
rect 230 194 231 195
rect 231 194 232 195
rect 232 194 233 195
rect 233 194 234 195
rect 360 194 361 195
rect 361 194 362 195
rect 362 194 363 195
rect 363 194 364 195
rect 364 194 365 195
rect 365 194 366 195
rect 366 194 367 195
rect 367 194 368 195
rect 368 194 369 195
rect 369 194 370 195
rect 370 194 371 195
rect 371 194 372 195
rect 372 194 373 195
rect 373 194 374 195
rect 374 194 375 195
rect 375 194 376 195
rect 376 194 377 195
rect 377 194 378 195
rect 378 194 379 195
rect 379 194 380 195
rect 380 194 381 195
rect 381 194 382 195
rect 382 194 383 195
rect 383 194 384 195
rect 384 194 385 195
rect 385 194 386 195
rect 386 194 387 195
rect 387 194 388 195
rect 388 194 389 195
rect 389 194 390 195
rect 390 194 391 195
rect 391 194 392 195
rect 392 194 393 195
rect 393 194 394 195
rect 394 194 395 195
rect 395 194 396 195
rect 396 194 397 195
rect 397 194 398 195
rect 398 194 399 195
rect 399 194 400 195
rect 400 194 401 195
rect 401 194 402 195
rect 402 194 403 195
rect 403 194 404 195
rect 404 194 405 195
rect 405 194 406 195
rect 406 194 407 195
rect 407 194 408 195
rect 433 194 434 195
rect 434 194 435 195
rect 435 194 436 195
rect 436 194 437 195
rect 437 194 438 195
rect 438 194 439 195
rect 439 194 440 195
rect 440 194 441 195
rect 441 194 442 195
rect 442 194 443 195
rect 443 194 444 195
rect 444 194 445 195
rect 514 194 515 195
rect 515 194 516 195
rect 516 194 517 195
rect 517 194 518 195
rect 518 194 519 195
rect 519 194 520 195
rect 520 194 521 195
rect 521 194 522 195
rect 522 194 523 195
rect 523 194 524 195
rect 524 194 525 195
rect 525 194 526 195
rect 526 194 527 195
rect 527 194 528 195
rect 94 193 95 194
rect 95 193 96 194
rect 96 193 97 194
rect 97 193 98 194
rect 98 193 99 194
rect 99 193 100 194
rect 100 193 101 194
rect 101 193 102 194
rect 102 193 103 194
rect 103 193 104 194
rect 165 193 166 194
rect 166 193 167 194
rect 167 193 168 194
rect 169 193 170 194
rect 170 193 171 194
rect 171 193 172 194
rect 172 193 173 194
rect 173 193 174 194
rect 174 193 175 194
rect 175 193 176 194
rect 176 193 177 194
rect 177 193 178 194
rect 178 193 179 194
rect 179 193 180 194
rect 180 193 181 194
rect 203 193 204 194
rect 204 193 205 194
rect 205 193 206 194
rect 206 193 207 194
rect 208 193 209 194
rect 209 193 210 194
rect 210 193 211 194
rect 211 193 212 194
rect 212 193 213 194
rect 214 193 215 194
rect 215 193 216 194
rect 216 193 217 194
rect 217 193 218 194
rect 218 193 219 194
rect 220 193 221 194
rect 221 193 222 194
rect 222 193 223 194
rect 223 193 224 194
rect 224 193 225 194
rect 225 193 226 194
rect 226 193 227 194
rect 227 193 228 194
rect 228 193 229 194
rect 229 193 230 194
rect 230 193 231 194
rect 231 193 232 194
rect 232 193 233 194
rect 233 193 234 194
rect 360 193 361 194
rect 361 193 362 194
rect 362 193 363 194
rect 363 193 364 194
rect 364 193 365 194
rect 365 193 366 194
rect 366 193 367 194
rect 367 193 368 194
rect 368 193 369 194
rect 369 193 370 194
rect 370 193 371 194
rect 371 193 372 194
rect 372 193 373 194
rect 373 193 374 194
rect 374 193 375 194
rect 375 193 376 194
rect 376 193 377 194
rect 377 193 378 194
rect 378 193 379 194
rect 379 193 380 194
rect 380 193 381 194
rect 381 193 382 194
rect 382 193 383 194
rect 383 193 384 194
rect 384 193 385 194
rect 385 193 386 194
rect 386 193 387 194
rect 387 193 388 194
rect 388 193 389 194
rect 389 193 390 194
rect 390 193 391 194
rect 391 193 392 194
rect 392 193 393 194
rect 393 193 394 194
rect 394 193 395 194
rect 395 193 396 194
rect 396 193 397 194
rect 397 193 398 194
rect 398 193 399 194
rect 399 193 400 194
rect 400 193 401 194
rect 401 193 402 194
rect 402 193 403 194
rect 403 193 404 194
rect 404 193 405 194
rect 405 193 406 194
rect 406 193 407 194
rect 407 193 408 194
rect 433 193 434 194
rect 434 193 435 194
rect 435 193 436 194
rect 436 193 437 194
rect 437 193 438 194
rect 438 193 439 194
rect 439 193 440 194
rect 440 193 441 194
rect 441 193 442 194
rect 442 193 443 194
rect 443 193 444 194
rect 444 193 445 194
rect 514 193 515 194
rect 515 193 516 194
rect 516 193 517 194
rect 517 193 518 194
rect 518 193 519 194
rect 519 193 520 194
rect 520 193 521 194
rect 521 193 522 194
rect 522 193 523 194
rect 523 193 524 194
rect 524 193 525 194
rect 525 193 526 194
rect 526 193 527 194
rect 527 193 528 194
rect 96 192 97 193
rect 97 192 98 193
rect 98 192 99 193
rect 99 192 100 193
rect 100 192 101 193
rect 101 192 102 193
rect 102 192 103 193
rect 103 192 104 193
rect 221 192 222 193
rect 222 192 223 193
rect 223 192 224 193
rect 224 192 225 193
rect 225 192 226 193
rect 226 192 227 193
rect 227 192 228 193
rect 228 192 229 193
rect 229 192 230 193
rect 230 192 231 193
rect 231 192 232 193
rect 232 192 233 193
rect 233 192 234 193
rect 362 192 363 193
rect 363 192 364 193
rect 364 192 365 193
rect 365 192 366 193
rect 366 192 367 193
rect 367 192 368 193
rect 368 192 369 193
rect 369 192 370 193
rect 370 192 371 193
rect 371 192 372 193
rect 372 192 373 193
rect 373 192 374 193
rect 374 192 375 193
rect 375 192 376 193
rect 376 192 377 193
rect 377 192 378 193
rect 378 192 379 193
rect 379 192 380 193
rect 380 192 381 193
rect 381 192 382 193
rect 382 192 383 193
rect 383 192 384 193
rect 384 192 385 193
rect 385 192 386 193
rect 386 192 387 193
rect 387 192 388 193
rect 388 192 389 193
rect 389 192 390 193
rect 390 192 391 193
rect 391 192 392 193
rect 392 192 393 193
rect 393 192 394 193
rect 394 192 395 193
rect 395 192 396 193
rect 396 192 397 193
rect 397 192 398 193
rect 398 192 399 193
rect 399 192 400 193
rect 400 192 401 193
rect 401 192 402 193
rect 402 192 403 193
rect 403 192 404 193
rect 404 192 405 193
rect 405 192 406 193
rect 406 192 407 193
rect 407 192 408 193
rect 435 192 436 193
rect 436 192 437 193
rect 437 192 438 193
rect 438 192 439 193
rect 439 192 440 193
rect 440 192 441 193
rect 441 192 442 193
rect 442 192 443 193
rect 443 192 444 193
rect 444 192 445 193
rect 514 192 515 193
rect 515 192 516 193
rect 516 192 517 193
rect 517 192 518 193
rect 518 192 519 193
rect 519 192 520 193
rect 520 192 521 193
rect 521 192 522 193
rect 522 192 523 193
rect 523 192 524 193
rect 524 192 525 193
rect 525 192 526 193
rect 526 192 527 193
rect 527 192 528 193
rect 96 191 97 192
rect 97 191 98 192
rect 98 191 99 192
rect 99 191 100 192
rect 100 191 101 192
rect 101 191 102 192
rect 102 191 103 192
rect 103 191 104 192
rect 104 191 105 192
rect 105 191 106 192
rect 221 191 222 192
rect 222 191 223 192
rect 223 191 224 192
rect 224 191 225 192
rect 225 191 226 192
rect 226 191 227 192
rect 227 191 228 192
rect 228 191 229 192
rect 229 191 230 192
rect 230 191 231 192
rect 231 191 232 192
rect 232 191 233 192
rect 233 191 234 192
rect 362 191 363 192
rect 363 191 364 192
rect 364 191 365 192
rect 365 191 366 192
rect 366 191 367 192
rect 367 191 368 192
rect 368 191 369 192
rect 369 191 370 192
rect 370 191 371 192
rect 371 191 372 192
rect 372 191 373 192
rect 373 191 374 192
rect 374 191 375 192
rect 375 191 376 192
rect 376 191 377 192
rect 377 191 378 192
rect 378 191 379 192
rect 379 191 380 192
rect 380 191 381 192
rect 381 191 382 192
rect 382 191 383 192
rect 383 191 384 192
rect 384 191 385 192
rect 385 191 386 192
rect 386 191 387 192
rect 387 191 388 192
rect 388 191 389 192
rect 389 191 390 192
rect 390 191 391 192
rect 391 191 392 192
rect 392 191 393 192
rect 393 191 394 192
rect 394 191 395 192
rect 395 191 396 192
rect 396 191 397 192
rect 397 191 398 192
rect 398 191 399 192
rect 399 191 400 192
rect 400 191 401 192
rect 401 191 402 192
rect 402 191 403 192
rect 403 191 404 192
rect 404 191 405 192
rect 405 191 406 192
rect 406 191 407 192
rect 407 191 408 192
rect 435 191 436 192
rect 436 191 437 192
rect 437 191 438 192
rect 438 191 439 192
rect 439 191 440 192
rect 440 191 441 192
rect 441 191 442 192
rect 442 191 443 192
rect 443 191 444 192
rect 444 191 445 192
rect 514 191 515 192
rect 515 191 516 192
rect 516 191 517 192
rect 517 191 518 192
rect 518 191 519 192
rect 519 191 520 192
rect 520 191 521 192
rect 521 191 522 192
rect 522 191 523 192
rect 523 191 524 192
rect 524 191 525 192
rect 525 191 526 192
rect 526 191 527 192
rect 527 191 528 192
rect 96 190 97 191
rect 97 190 98 191
rect 98 190 99 191
rect 99 190 100 191
rect 100 190 101 191
rect 101 190 102 191
rect 102 190 103 191
rect 103 190 104 191
rect 104 190 105 191
rect 105 190 106 191
rect 221 190 222 191
rect 222 190 223 191
rect 223 190 224 191
rect 224 190 225 191
rect 225 190 226 191
rect 226 190 227 191
rect 227 190 228 191
rect 228 190 229 191
rect 229 190 230 191
rect 230 190 231 191
rect 231 190 232 191
rect 232 190 233 191
rect 233 190 234 191
rect 364 190 365 191
rect 365 190 366 191
rect 366 190 367 191
rect 367 190 368 191
rect 368 190 369 191
rect 369 190 370 191
rect 370 190 371 191
rect 371 190 372 191
rect 372 190 373 191
rect 373 190 374 191
rect 374 190 375 191
rect 375 190 376 191
rect 376 190 377 191
rect 377 190 378 191
rect 399 190 400 191
rect 400 190 401 191
rect 401 190 402 191
rect 402 190 403 191
rect 403 190 404 191
rect 404 190 405 191
rect 405 190 406 191
rect 406 190 407 191
rect 407 190 408 191
rect 435 190 436 191
rect 436 190 437 191
rect 437 190 438 191
rect 438 190 439 191
rect 439 190 440 191
rect 440 190 441 191
rect 441 190 442 191
rect 442 190 443 191
rect 443 190 444 191
rect 444 190 445 191
rect 514 190 515 191
rect 515 190 516 191
rect 516 190 517 191
rect 517 190 518 191
rect 518 190 519 191
rect 519 190 520 191
rect 520 190 521 191
rect 521 190 522 191
rect 522 190 523 191
rect 523 190 524 191
rect 524 190 525 191
rect 525 190 526 191
rect 96 189 97 190
rect 97 189 98 190
rect 98 189 99 190
rect 99 189 100 190
rect 100 189 101 190
rect 101 189 102 190
rect 102 189 103 190
rect 103 189 104 190
rect 104 189 105 190
rect 105 189 106 190
rect 220 189 221 190
rect 221 189 222 190
rect 222 189 223 190
rect 223 189 224 190
rect 224 189 225 190
rect 225 189 226 190
rect 226 189 227 190
rect 227 189 228 190
rect 228 189 229 190
rect 229 189 230 190
rect 230 189 231 190
rect 231 189 232 190
rect 232 189 233 190
rect 233 189 234 190
rect 234 189 235 190
rect 235 189 236 190
rect 289 189 290 190
rect 290 189 291 190
rect 291 189 292 190
rect 292 189 293 190
rect 293 189 294 190
rect 364 189 365 190
rect 365 189 366 190
rect 366 189 367 190
rect 367 189 368 190
rect 368 189 369 190
rect 369 189 370 190
rect 370 189 371 190
rect 371 189 372 190
rect 372 189 373 190
rect 373 189 374 190
rect 374 189 375 190
rect 375 189 376 190
rect 376 189 377 190
rect 377 189 378 190
rect 399 189 400 190
rect 400 189 401 190
rect 401 189 402 190
rect 402 189 403 190
rect 403 189 404 190
rect 404 189 405 190
rect 405 189 406 190
rect 406 189 407 190
rect 407 189 408 190
rect 433 189 434 190
rect 434 189 435 190
rect 435 189 436 190
rect 436 189 437 190
rect 437 189 438 190
rect 438 189 439 190
rect 439 189 440 190
rect 440 189 441 190
rect 441 189 442 190
rect 442 189 443 190
rect 443 189 444 190
rect 444 189 445 190
rect 512 189 513 190
rect 513 189 514 190
rect 514 189 515 190
rect 515 189 516 190
rect 516 189 517 190
rect 517 189 518 190
rect 518 189 519 190
rect 519 189 520 190
rect 520 189 521 190
rect 521 189 522 190
rect 522 189 523 190
rect 523 189 524 190
rect 524 189 525 190
rect 525 189 526 190
rect 96 188 97 189
rect 97 188 98 189
rect 98 188 99 189
rect 99 188 100 189
rect 100 188 101 189
rect 101 188 102 189
rect 102 188 103 189
rect 103 188 104 189
rect 104 188 105 189
rect 105 188 106 189
rect 220 188 221 189
rect 221 188 222 189
rect 222 188 223 189
rect 223 188 224 189
rect 224 188 225 189
rect 225 188 226 189
rect 226 188 227 189
rect 227 188 228 189
rect 228 188 229 189
rect 229 188 230 189
rect 230 188 231 189
rect 231 188 232 189
rect 232 188 233 189
rect 233 188 234 189
rect 234 188 235 189
rect 235 188 236 189
rect 289 188 290 189
rect 290 188 291 189
rect 291 188 292 189
rect 292 188 293 189
rect 293 188 294 189
rect 366 188 367 189
rect 367 188 368 189
rect 368 188 369 189
rect 369 188 370 189
rect 370 188 371 189
rect 371 188 372 189
rect 372 188 373 189
rect 373 188 374 189
rect 374 188 375 189
rect 375 188 376 189
rect 376 188 377 189
rect 377 188 378 189
rect 401 188 402 189
rect 402 188 403 189
rect 403 188 404 189
rect 404 188 405 189
rect 405 188 406 189
rect 406 188 407 189
rect 407 188 408 189
rect 433 188 434 189
rect 434 188 435 189
rect 435 188 436 189
rect 436 188 437 189
rect 437 188 438 189
rect 438 188 439 189
rect 439 188 440 189
rect 440 188 441 189
rect 441 188 442 189
rect 442 188 443 189
rect 443 188 444 189
rect 444 188 445 189
rect 512 188 513 189
rect 513 188 514 189
rect 514 188 515 189
rect 515 188 516 189
rect 516 188 517 189
rect 517 188 518 189
rect 518 188 519 189
rect 519 188 520 189
rect 520 188 521 189
rect 521 188 522 189
rect 522 188 523 189
rect 523 188 524 189
rect 524 188 525 189
rect 525 188 526 189
rect 96 187 97 188
rect 97 187 98 188
rect 98 187 99 188
rect 99 187 100 188
rect 100 187 101 188
rect 101 187 102 188
rect 102 187 103 188
rect 103 187 104 188
rect 104 187 105 188
rect 105 187 106 188
rect 220 187 221 188
rect 221 187 222 188
rect 222 187 223 188
rect 223 187 224 188
rect 224 187 225 188
rect 225 187 226 188
rect 226 187 227 188
rect 227 187 228 188
rect 228 187 229 188
rect 229 187 230 188
rect 230 187 231 188
rect 231 187 232 188
rect 232 187 233 188
rect 233 187 234 188
rect 234 187 235 188
rect 235 187 236 188
rect 289 187 290 188
rect 290 187 291 188
rect 291 187 292 188
rect 292 187 293 188
rect 293 187 294 188
rect 366 187 367 188
rect 367 187 368 188
rect 368 187 369 188
rect 369 187 370 188
rect 370 187 371 188
rect 371 187 372 188
rect 372 187 373 188
rect 373 187 374 188
rect 374 187 375 188
rect 375 187 376 188
rect 376 187 377 188
rect 377 187 378 188
rect 378 187 379 188
rect 379 187 380 188
rect 401 187 402 188
rect 402 187 403 188
rect 403 187 404 188
rect 404 187 405 188
rect 405 187 406 188
rect 406 187 407 188
rect 407 187 408 188
rect 433 187 434 188
rect 434 187 435 188
rect 435 187 436 188
rect 436 187 437 188
rect 437 187 438 188
rect 438 187 439 188
rect 439 187 440 188
rect 440 187 441 188
rect 441 187 442 188
rect 442 187 443 188
rect 443 187 444 188
rect 444 187 445 188
rect 510 187 511 188
rect 511 187 512 188
rect 512 187 513 188
rect 513 187 514 188
rect 514 187 515 188
rect 515 187 516 188
rect 516 187 517 188
rect 517 187 518 188
rect 518 187 519 188
rect 519 187 520 188
rect 520 187 521 188
rect 521 187 522 188
rect 522 187 523 188
rect 523 187 524 188
rect 524 187 525 188
rect 525 187 526 188
rect 98 186 99 187
rect 99 186 100 187
rect 100 186 101 187
rect 101 186 102 187
rect 102 186 103 187
rect 103 186 104 187
rect 104 186 105 187
rect 105 186 106 187
rect 220 186 221 187
rect 221 186 222 187
rect 222 186 223 187
rect 223 186 224 187
rect 224 186 225 187
rect 225 186 226 187
rect 226 186 227 187
rect 227 186 228 187
rect 228 186 229 187
rect 229 186 230 187
rect 230 186 231 187
rect 231 186 232 187
rect 232 186 233 187
rect 233 186 234 187
rect 234 186 235 187
rect 235 186 236 187
rect 289 186 290 187
rect 290 186 291 187
rect 291 186 292 187
rect 292 186 293 187
rect 293 186 294 187
rect 366 186 367 187
rect 367 186 368 187
rect 368 186 369 187
rect 369 186 370 187
rect 370 186 371 187
rect 371 186 372 187
rect 372 186 373 187
rect 373 186 374 187
rect 374 186 375 187
rect 375 186 376 187
rect 376 186 377 187
rect 377 186 378 187
rect 378 186 379 187
rect 379 186 380 187
rect 403 186 404 187
rect 404 186 405 187
rect 405 186 406 187
rect 406 186 407 187
rect 407 186 408 187
rect 435 186 436 187
rect 436 186 437 187
rect 437 186 438 187
rect 438 186 439 187
rect 439 186 440 187
rect 440 186 441 187
rect 441 186 442 187
rect 442 186 443 187
rect 443 186 444 187
rect 444 186 445 187
rect 510 186 511 187
rect 511 186 512 187
rect 512 186 513 187
rect 513 186 514 187
rect 514 186 515 187
rect 515 186 516 187
rect 516 186 517 187
rect 517 186 518 187
rect 518 186 519 187
rect 519 186 520 187
rect 520 186 521 187
rect 521 186 522 187
rect 522 186 523 187
rect 523 186 524 187
rect 98 185 99 186
rect 99 185 100 186
rect 100 185 101 186
rect 101 185 102 186
rect 102 185 103 186
rect 103 185 104 186
rect 104 185 105 186
rect 105 185 106 186
rect 106 185 107 186
rect 107 185 108 186
rect 220 185 221 186
rect 221 185 222 186
rect 222 185 223 186
rect 223 185 224 186
rect 224 185 225 186
rect 225 185 226 186
rect 226 185 227 186
rect 227 185 228 186
rect 228 185 229 186
rect 229 185 230 186
rect 230 185 231 186
rect 231 185 232 186
rect 232 185 233 186
rect 233 185 234 186
rect 234 185 235 186
rect 235 185 236 186
rect 236 185 237 186
rect 287 185 288 186
rect 288 185 289 186
rect 289 185 290 186
rect 290 185 291 186
rect 291 185 292 186
rect 292 185 293 186
rect 293 185 294 186
rect 294 185 295 186
rect 366 185 367 186
rect 367 185 368 186
rect 368 185 369 186
rect 369 185 370 186
rect 370 185 371 186
rect 371 185 372 186
rect 372 185 373 186
rect 373 185 374 186
rect 374 185 375 186
rect 375 185 376 186
rect 376 185 377 186
rect 377 185 378 186
rect 378 185 379 186
rect 379 185 380 186
rect 380 185 381 186
rect 381 185 382 186
rect 403 185 404 186
rect 404 185 405 186
rect 405 185 406 186
rect 406 185 407 186
rect 407 185 408 186
rect 435 185 436 186
rect 436 185 437 186
rect 437 185 438 186
rect 438 185 439 186
rect 439 185 440 186
rect 440 185 441 186
rect 441 185 442 186
rect 442 185 443 186
rect 443 185 444 186
rect 444 185 445 186
rect 510 185 511 186
rect 511 185 512 186
rect 512 185 513 186
rect 513 185 514 186
rect 514 185 515 186
rect 515 185 516 186
rect 516 185 517 186
rect 517 185 518 186
rect 518 185 519 186
rect 519 185 520 186
rect 520 185 521 186
rect 521 185 522 186
rect 522 185 523 186
rect 523 185 524 186
rect 98 184 99 185
rect 99 184 100 185
rect 100 184 101 185
rect 101 184 102 185
rect 102 184 103 185
rect 103 184 104 185
rect 104 184 105 185
rect 105 184 106 185
rect 106 184 107 185
rect 107 184 108 185
rect 220 184 221 185
rect 221 184 222 185
rect 222 184 223 185
rect 223 184 224 185
rect 225 184 226 185
rect 226 184 227 185
rect 227 184 228 185
rect 228 184 229 185
rect 229 184 230 185
rect 230 184 231 185
rect 231 184 232 185
rect 232 184 233 185
rect 233 184 234 185
rect 234 184 235 185
rect 235 184 236 185
rect 236 184 237 185
rect 287 184 288 185
rect 288 184 289 185
rect 289 184 290 185
rect 290 184 291 185
rect 291 184 292 185
rect 292 184 293 185
rect 293 184 294 185
rect 294 184 295 185
rect 368 184 369 185
rect 369 184 370 185
rect 370 184 371 185
rect 371 184 372 185
rect 372 184 373 185
rect 373 184 374 185
rect 374 184 375 185
rect 375 184 376 185
rect 376 184 377 185
rect 377 184 378 185
rect 378 184 379 185
rect 379 184 380 185
rect 380 184 381 185
rect 381 184 382 185
rect 405 184 406 185
rect 406 184 407 185
rect 407 184 408 185
rect 435 184 436 185
rect 436 184 437 185
rect 437 184 438 185
rect 438 184 439 185
rect 439 184 440 185
rect 440 184 441 185
rect 441 184 442 185
rect 442 184 443 185
rect 443 184 444 185
rect 444 184 445 185
rect 510 184 511 185
rect 511 184 512 185
rect 512 184 513 185
rect 513 184 514 185
rect 514 184 515 185
rect 515 184 516 185
rect 516 184 517 185
rect 517 184 518 185
rect 518 184 519 185
rect 519 184 520 185
rect 520 184 521 185
rect 521 184 522 185
rect 522 184 523 185
rect 523 184 524 185
rect 98 183 99 184
rect 99 183 100 184
rect 100 183 101 184
rect 101 183 102 184
rect 102 183 103 184
rect 103 183 104 184
rect 104 183 105 184
rect 105 183 106 184
rect 106 183 107 184
rect 107 183 108 184
rect 220 183 221 184
rect 221 183 222 184
rect 222 183 223 184
rect 223 183 224 184
rect 225 183 226 184
rect 226 183 227 184
rect 227 183 228 184
rect 228 183 229 184
rect 229 183 230 184
rect 230 183 231 184
rect 231 183 232 184
rect 232 183 233 184
rect 233 183 234 184
rect 234 183 235 184
rect 235 183 236 184
rect 236 183 237 184
rect 287 183 288 184
rect 288 183 289 184
rect 289 183 290 184
rect 290 183 291 184
rect 291 183 292 184
rect 292 183 293 184
rect 293 183 294 184
rect 294 183 295 184
rect 368 183 369 184
rect 369 183 370 184
rect 370 183 371 184
rect 371 183 372 184
rect 372 183 373 184
rect 373 183 374 184
rect 374 183 375 184
rect 375 183 376 184
rect 376 183 377 184
rect 377 183 378 184
rect 378 183 379 184
rect 379 183 380 184
rect 380 183 381 184
rect 381 183 382 184
rect 382 183 383 184
rect 383 183 384 184
rect 405 183 406 184
rect 406 183 407 184
rect 407 183 408 184
rect 433 183 434 184
rect 434 183 435 184
rect 435 183 436 184
rect 436 183 437 184
rect 437 183 438 184
rect 438 183 439 184
rect 439 183 440 184
rect 440 183 441 184
rect 441 183 442 184
rect 442 183 443 184
rect 443 183 444 184
rect 444 183 445 184
rect 508 183 509 184
rect 509 183 510 184
rect 510 183 511 184
rect 511 183 512 184
rect 512 183 513 184
rect 513 183 514 184
rect 514 183 515 184
rect 515 183 516 184
rect 516 183 517 184
rect 517 183 518 184
rect 518 183 519 184
rect 519 183 520 184
rect 520 183 521 184
rect 521 183 522 184
rect 522 183 523 184
rect 523 183 524 184
rect 98 182 99 183
rect 99 182 100 183
rect 100 182 101 183
rect 101 182 102 183
rect 102 182 103 183
rect 103 182 104 183
rect 104 182 105 183
rect 105 182 106 183
rect 106 182 107 183
rect 107 182 108 183
rect 220 182 221 183
rect 221 182 222 183
rect 222 182 223 183
rect 223 182 224 183
rect 227 182 228 183
rect 228 182 229 183
rect 229 182 230 183
rect 230 182 231 183
rect 231 182 232 183
rect 232 182 233 183
rect 233 182 234 183
rect 234 182 235 183
rect 235 182 236 183
rect 236 182 237 183
rect 287 182 288 183
rect 288 182 289 183
rect 289 182 290 183
rect 290 182 291 183
rect 291 182 292 183
rect 292 182 293 183
rect 293 182 294 183
rect 294 182 295 183
rect 369 182 370 183
rect 370 182 371 183
rect 371 182 372 183
rect 372 182 373 183
rect 373 182 374 183
rect 374 182 375 183
rect 375 182 376 183
rect 376 182 377 183
rect 377 182 378 183
rect 378 182 379 183
rect 379 182 380 183
rect 380 182 381 183
rect 381 182 382 183
rect 382 182 383 183
rect 383 182 384 183
rect 405 182 406 183
rect 406 182 407 183
rect 407 182 408 183
rect 433 182 434 183
rect 434 182 435 183
rect 435 182 436 183
rect 436 182 437 183
rect 437 182 438 183
rect 438 182 439 183
rect 439 182 440 183
rect 440 182 441 183
rect 441 182 442 183
rect 442 182 443 183
rect 443 182 444 183
rect 444 182 445 183
rect 508 182 509 183
rect 509 182 510 183
rect 510 182 511 183
rect 511 182 512 183
rect 512 182 513 183
rect 513 182 514 183
rect 514 182 515 183
rect 515 182 516 183
rect 516 182 517 183
rect 517 182 518 183
rect 518 182 519 183
rect 519 182 520 183
rect 520 182 521 183
rect 521 182 522 183
rect 522 182 523 183
rect 523 182 524 183
rect 98 181 99 182
rect 99 181 100 182
rect 100 181 101 182
rect 101 181 102 182
rect 102 181 103 182
rect 103 181 104 182
rect 104 181 105 182
rect 105 181 106 182
rect 106 181 107 182
rect 107 181 108 182
rect 218 181 219 182
rect 219 181 220 182
rect 220 181 221 182
rect 221 181 222 182
rect 222 181 223 182
rect 223 181 224 182
rect 227 181 228 182
rect 228 181 229 182
rect 229 181 230 182
rect 230 181 231 182
rect 231 181 232 182
rect 232 181 233 182
rect 233 181 234 182
rect 234 181 235 182
rect 235 181 236 182
rect 236 181 237 182
rect 237 181 238 182
rect 238 181 239 182
rect 287 181 288 182
rect 288 181 289 182
rect 289 181 290 182
rect 290 181 291 182
rect 291 181 292 182
rect 292 181 293 182
rect 293 181 294 182
rect 294 181 295 182
rect 369 181 370 182
rect 370 181 371 182
rect 371 181 372 182
rect 372 181 373 182
rect 373 181 374 182
rect 374 181 375 182
rect 375 181 376 182
rect 376 181 377 182
rect 377 181 378 182
rect 378 181 379 182
rect 379 181 380 182
rect 380 181 381 182
rect 381 181 382 182
rect 382 181 383 182
rect 383 181 384 182
rect 405 181 406 182
rect 406 181 407 182
rect 407 181 408 182
rect 433 181 434 182
rect 434 181 435 182
rect 435 181 436 182
rect 436 181 437 182
rect 437 181 438 182
rect 438 181 439 182
rect 439 181 440 182
rect 440 181 441 182
rect 441 181 442 182
rect 442 181 443 182
rect 443 181 444 182
rect 444 181 445 182
rect 508 181 509 182
rect 509 181 510 182
rect 510 181 511 182
rect 511 181 512 182
rect 512 181 513 182
rect 513 181 514 182
rect 514 181 515 182
rect 515 181 516 182
rect 516 181 517 182
rect 517 181 518 182
rect 518 181 519 182
rect 519 181 520 182
rect 520 181 521 182
rect 521 181 522 182
rect 522 181 523 182
rect 523 181 524 182
rect 100 180 101 181
rect 101 180 102 181
rect 102 180 103 181
rect 103 180 104 181
rect 104 180 105 181
rect 105 180 106 181
rect 106 180 107 181
rect 107 180 108 181
rect 218 180 219 181
rect 219 180 220 181
rect 220 180 221 181
rect 221 180 222 181
rect 222 180 223 181
rect 223 180 224 181
rect 227 180 228 181
rect 228 180 229 181
rect 229 180 230 181
rect 230 180 231 181
rect 231 180 232 181
rect 232 180 233 181
rect 233 180 234 181
rect 234 180 235 181
rect 235 180 236 181
rect 236 180 237 181
rect 237 180 238 181
rect 238 180 239 181
rect 287 180 288 181
rect 288 180 289 181
rect 289 180 290 181
rect 290 180 291 181
rect 291 180 292 181
rect 292 180 293 181
rect 293 180 294 181
rect 294 180 295 181
rect 371 180 372 181
rect 372 180 373 181
rect 373 180 374 181
rect 374 180 375 181
rect 375 180 376 181
rect 376 180 377 181
rect 377 180 378 181
rect 378 180 379 181
rect 379 180 380 181
rect 380 180 381 181
rect 381 180 382 181
rect 382 180 383 181
rect 383 180 384 181
rect 435 180 436 181
rect 436 180 437 181
rect 437 180 438 181
rect 438 180 439 181
rect 439 180 440 181
rect 440 180 441 181
rect 441 180 442 181
rect 442 180 443 181
rect 443 180 444 181
rect 444 180 445 181
rect 508 180 509 181
rect 509 180 510 181
rect 510 180 511 181
rect 511 180 512 181
rect 512 180 513 181
rect 513 180 514 181
rect 514 180 515 181
rect 515 180 516 181
rect 516 180 517 181
rect 517 180 518 181
rect 518 180 519 181
rect 519 180 520 181
rect 520 180 521 181
rect 521 180 522 181
rect 100 179 101 180
rect 101 179 102 180
rect 102 179 103 180
rect 103 179 104 180
rect 104 179 105 180
rect 105 179 106 180
rect 106 179 107 180
rect 107 179 108 180
rect 218 179 219 180
rect 219 179 220 180
rect 220 179 221 180
rect 221 179 222 180
rect 222 179 223 180
rect 223 179 224 180
rect 227 179 228 180
rect 228 179 229 180
rect 229 179 230 180
rect 230 179 231 180
rect 231 179 232 180
rect 232 179 233 180
rect 233 179 234 180
rect 234 179 235 180
rect 235 179 236 180
rect 236 179 237 180
rect 237 179 238 180
rect 238 179 239 180
rect 287 179 288 180
rect 288 179 289 180
rect 289 179 290 180
rect 290 179 291 180
rect 291 179 292 180
rect 292 179 293 180
rect 293 179 294 180
rect 294 179 295 180
rect 371 179 372 180
rect 372 179 373 180
rect 373 179 374 180
rect 374 179 375 180
rect 375 179 376 180
rect 376 179 377 180
rect 377 179 378 180
rect 378 179 379 180
rect 379 179 380 180
rect 380 179 381 180
rect 381 179 382 180
rect 382 179 383 180
rect 383 179 384 180
rect 435 179 436 180
rect 436 179 437 180
rect 437 179 438 180
rect 438 179 439 180
rect 439 179 440 180
rect 440 179 441 180
rect 441 179 442 180
rect 442 179 443 180
rect 443 179 444 180
rect 444 179 445 180
rect 508 179 509 180
rect 509 179 510 180
rect 510 179 511 180
rect 511 179 512 180
rect 512 179 513 180
rect 513 179 514 180
rect 514 179 515 180
rect 515 179 516 180
rect 516 179 517 180
rect 517 179 518 180
rect 518 179 519 180
rect 519 179 520 180
rect 520 179 521 180
rect 521 179 522 180
rect 100 178 101 179
rect 101 178 102 179
rect 102 178 103 179
rect 103 178 104 179
rect 104 178 105 179
rect 105 178 106 179
rect 106 178 107 179
rect 107 178 108 179
rect 108 178 109 179
rect 109 178 110 179
rect 216 178 217 179
rect 217 178 218 179
rect 218 178 219 179
rect 219 178 220 179
rect 220 178 221 179
rect 221 178 222 179
rect 222 178 223 179
rect 223 178 224 179
rect 227 178 228 179
rect 228 178 229 179
rect 229 178 230 179
rect 230 178 231 179
rect 231 178 232 179
rect 232 178 233 179
rect 233 178 234 179
rect 234 178 235 179
rect 235 178 236 179
rect 236 178 237 179
rect 237 178 238 179
rect 238 178 239 179
rect 285 178 286 179
rect 286 178 287 179
rect 287 178 288 179
rect 288 178 289 179
rect 289 178 290 179
rect 290 178 291 179
rect 291 178 292 179
rect 292 178 293 179
rect 293 178 294 179
rect 294 178 295 179
rect 295 178 296 179
rect 296 178 297 179
rect 371 178 372 179
rect 372 178 373 179
rect 373 178 374 179
rect 374 178 375 179
rect 375 178 376 179
rect 376 178 377 179
rect 377 178 378 179
rect 378 178 379 179
rect 379 178 380 179
rect 380 178 381 179
rect 381 178 382 179
rect 382 178 383 179
rect 383 178 384 179
rect 384 178 385 179
rect 433 178 434 179
rect 434 178 435 179
rect 435 178 436 179
rect 436 178 437 179
rect 437 178 438 179
rect 438 178 439 179
rect 439 178 440 179
rect 440 178 441 179
rect 441 178 442 179
rect 442 178 443 179
rect 443 178 444 179
rect 444 178 445 179
rect 506 178 507 179
rect 507 178 508 179
rect 508 178 509 179
rect 509 178 510 179
rect 510 178 511 179
rect 511 178 512 179
rect 512 178 513 179
rect 513 178 514 179
rect 514 178 515 179
rect 515 178 516 179
rect 516 178 517 179
rect 517 178 518 179
rect 518 178 519 179
rect 519 178 520 179
rect 520 178 521 179
rect 521 178 522 179
rect 100 177 101 178
rect 101 177 102 178
rect 102 177 103 178
rect 103 177 104 178
rect 104 177 105 178
rect 105 177 106 178
rect 106 177 107 178
rect 107 177 108 178
rect 108 177 109 178
rect 109 177 110 178
rect 216 177 217 178
rect 217 177 218 178
rect 218 177 219 178
rect 219 177 220 178
rect 220 177 221 178
rect 221 177 222 178
rect 227 177 228 178
rect 228 177 229 178
rect 229 177 230 178
rect 230 177 231 178
rect 231 177 232 178
rect 232 177 233 178
rect 233 177 234 178
rect 234 177 235 178
rect 235 177 236 178
rect 236 177 237 178
rect 237 177 238 178
rect 238 177 239 178
rect 285 177 286 178
rect 286 177 287 178
rect 287 177 288 178
rect 288 177 289 178
rect 289 177 290 178
rect 290 177 291 178
rect 291 177 292 178
rect 292 177 293 178
rect 293 177 294 178
rect 294 177 295 178
rect 295 177 296 178
rect 296 177 297 178
rect 371 177 372 178
rect 372 177 373 178
rect 373 177 374 178
rect 374 177 375 178
rect 375 177 376 178
rect 376 177 377 178
rect 377 177 378 178
rect 378 177 379 178
rect 379 177 380 178
rect 380 177 381 178
rect 381 177 382 178
rect 382 177 383 178
rect 383 177 384 178
rect 384 177 385 178
rect 433 177 434 178
rect 434 177 435 178
rect 435 177 436 178
rect 436 177 437 178
rect 437 177 438 178
rect 438 177 439 178
rect 439 177 440 178
rect 440 177 441 178
rect 441 177 442 178
rect 442 177 443 178
rect 443 177 444 178
rect 444 177 445 178
rect 506 177 507 178
rect 507 177 508 178
rect 508 177 509 178
rect 509 177 510 178
rect 510 177 511 178
rect 511 177 512 178
rect 512 177 513 178
rect 513 177 514 178
rect 514 177 515 178
rect 515 177 516 178
rect 516 177 517 178
rect 517 177 518 178
rect 518 177 519 178
rect 519 177 520 178
rect 520 177 521 178
rect 521 177 522 178
rect 100 176 101 177
rect 101 176 102 177
rect 102 176 103 177
rect 103 176 104 177
rect 104 176 105 177
rect 105 176 106 177
rect 106 176 107 177
rect 107 176 108 177
rect 108 176 109 177
rect 109 176 110 177
rect 216 176 217 177
rect 217 176 218 177
rect 218 176 219 177
rect 219 176 220 177
rect 220 176 221 177
rect 221 176 222 177
rect 227 176 228 177
rect 228 176 229 177
rect 229 176 230 177
rect 230 176 231 177
rect 231 176 232 177
rect 232 176 233 177
rect 233 176 234 177
rect 234 176 235 177
rect 235 176 236 177
rect 236 176 237 177
rect 237 176 238 177
rect 238 176 239 177
rect 285 176 286 177
rect 286 176 287 177
rect 287 176 288 177
rect 288 176 289 177
rect 289 176 290 177
rect 290 176 291 177
rect 291 176 292 177
rect 292 176 293 177
rect 293 176 294 177
rect 294 176 295 177
rect 295 176 296 177
rect 296 176 297 177
rect 328 176 329 177
rect 329 176 330 177
rect 330 176 331 177
rect 331 176 332 177
rect 332 176 333 177
rect 333 176 334 177
rect 334 176 335 177
rect 335 176 336 177
rect 336 176 337 177
rect 337 176 338 177
rect 338 176 339 177
rect 339 176 340 177
rect 340 176 341 177
rect 341 176 342 177
rect 342 176 343 177
rect 343 176 344 177
rect 344 176 345 177
rect 345 176 346 177
rect 346 176 347 177
rect 347 176 348 177
rect 348 176 349 177
rect 349 176 350 177
rect 351 176 352 177
rect 352 176 353 177
rect 353 176 354 177
rect 371 176 372 177
rect 372 176 373 177
rect 373 176 374 177
rect 374 176 375 177
rect 375 176 376 177
rect 376 176 377 177
rect 377 176 378 177
rect 378 176 379 177
rect 379 176 380 177
rect 380 176 381 177
rect 381 176 382 177
rect 382 176 383 177
rect 383 176 384 177
rect 384 176 385 177
rect 385 176 386 177
rect 386 176 387 177
rect 433 176 434 177
rect 434 176 435 177
rect 435 176 436 177
rect 436 176 437 177
rect 437 176 438 177
rect 438 176 439 177
rect 439 176 440 177
rect 440 176 441 177
rect 441 176 442 177
rect 442 176 443 177
rect 443 176 444 177
rect 444 176 445 177
rect 504 176 505 177
rect 505 176 506 177
rect 506 176 507 177
rect 507 176 508 177
rect 508 176 509 177
rect 509 176 510 177
rect 510 176 511 177
rect 511 176 512 177
rect 512 176 513 177
rect 513 176 514 177
rect 514 176 515 177
rect 515 176 516 177
rect 516 176 517 177
rect 517 176 518 177
rect 518 176 519 177
rect 519 176 520 177
rect 520 176 521 177
rect 521 176 522 177
rect 100 175 101 176
rect 101 175 102 176
rect 102 175 103 176
rect 103 175 104 176
rect 104 175 105 176
rect 105 175 106 176
rect 106 175 107 176
rect 107 175 108 176
rect 108 175 109 176
rect 109 175 110 176
rect 216 175 217 176
rect 217 175 218 176
rect 218 175 219 176
rect 219 175 220 176
rect 220 175 221 176
rect 221 175 222 176
rect 229 175 230 176
rect 230 175 231 176
rect 231 175 232 176
rect 232 175 233 176
rect 233 175 234 176
rect 234 175 235 176
rect 235 175 236 176
rect 236 175 237 176
rect 237 175 238 176
rect 238 175 239 176
rect 285 175 286 176
rect 286 175 287 176
rect 287 175 288 176
rect 288 175 289 176
rect 289 175 290 176
rect 290 175 291 176
rect 291 175 292 176
rect 292 175 293 176
rect 293 175 294 176
rect 294 175 295 176
rect 295 175 296 176
rect 296 175 297 176
rect 328 175 329 176
rect 329 175 330 176
rect 330 175 331 176
rect 331 175 332 176
rect 332 175 333 176
rect 333 175 334 176
rect 334 175 335 176
rect 335 175 336 176
rect 336 175 337 176
rect 337 175 338 176
rect 338 175 339 176
rect 339 175 340 176
rect 340 175 341 176
rect 341 175 342 176
rect 342 175 343 176
rect 343 175 344 176
rect 344 175 345 176
rect 345 175 346 176
rect 346 175 347 176
rect 347 175 348 176
rect 348 175 349 176
rect 349 175 350 176
rect 351 175 352 176
rect 352 175 353 176
rect 353 175 354 176
rect 373 175 374 176
rect 374 175 375 176
rect 375 175 376 176
rect 376 175 377 176
rect 377 175 378 176
rect 378 175 379 176
rect 379 175 380 176
rect 380 175 381 176
rect 381 175 382 176
rect 382 175 383 176
rect 383 175 384 176
rect 384 175 385 176
rect 385 175 386 176
rect 386 175 387 176
rect 435 175 436 176
rect 436 175 437 176
rect 437 175 438 176
rect 438 175 439 176
rect 439 175 440 176
rect 440 175 441 176
rect 441 175 442 176
rect 442 175 443 176
rect 443 175 444 176
rect 444 175 445 176
rect 504 175 505 176
rect 505 175 506 176
rect 506 175 507 176
rect 507 175 508 176
rect 508 175 509 176
rect 509 175 510 176
rect 510 175 511 176
rect 511 175 512 176
rect 512 175 513 176
rect 513 175 514 176
rect 514 175 515 176
rect 515 175 516 176
rect 516 175 517 176
rect 517 175 518 176
rect 518 175 519 176
rect 519 175 520 176
rect 100 174 101 175
rect 101 174 102 175
rect 102 174 103 175
rect 103 174 104 175
rect 104 174 105 175
rect 105 174 106 175
rect 106 174 107 175
rect 107 174 108 175
rect 108 174 109 175
rect 109 174 110 175
rect 216 174 217 175
rect 217 174 218 175
rect 218 174 219 175
rect 219 174 220 175
rect 220 174 221 175
rect 221 174 222 175
rect 229 174 230 175
rect 230 174 231 175
rect 231 174 232 175
rect 232 174 233 175
rect 233 174 234 175
rect 234 174 235 175
rect 235 174 236 175
rect 236 174 237 175
rect 237 174 238 175
rect 238 174 239 175
rect 239 174 240 175
rect 240 174 241 175
rect 285 174 286 175
rect 286 174 287 175
rect 287 174 288 175
rect 288 174 289 175
rect 289 174 290 175
rect 290 174 291 175
rect 291 174 292 175
rect 292 174 293 175
rect 293 174 294 175
rect 294 174 295 175
rect 295 174 296 175
rect 296 174 297 175
rect 297 174 298 175
rect 298 174 299 175
rect 328 174 329 175
rect 329 174 330 175
rect 330 174 331 175
rect 331 174 332 175
rect 332 174 333 175
rect 333 174 334 175
rect 334 174 335 175
rect 335 174 336 175
rect 336 174 337 175
rect 337 174 338 175
rect 338 174 339 175
rect 339 174 340 175
rect 340 174 341 175
rect 341 174 342 175
rect 342 174 343 175
rect 343 174 344 175
rect 344 174 345 175
rect 345 174 346 175
rect 346 174 347 175
rect 347 174 348 175
rect 348 174 349 175
rect 349 174 350 175
rect 350 174 351 175
rect 351 174 352 175
rect 352 174 353 175
rect 353 174 354 175
rect 373 174 374 175
rect 374 174 375 175
rect 375 174 376 175
rect 376 174 377 175
rect 377 174 378 175
rect 378 174 379 175
rect 379 174 380 175
rect 380 174 381 175
rect 381 174 382 175
rect 382 174 383 175
rect 383 174 384 175
rect 384 174 385 175
rect 385 174 386 175
rect 386 174 387 175
rect 387 174 388 175
rect 388 174 389 175
rect 435 174 436 175
rect 436 174 437 175
rect 437 174 438 175
rect 438 174 439 175
rect 439 174 440 175
rect 440 174 441 175
rect 441 174 442 175
rect 442 174 443 175
rect 443 174 444 175
rect 444 174 445 175
rect 504 174 505 175
rect 505 174 506 175
rect 506 174 507 175
rect 507 174 508 175
rect 508 174 509 175
rect 509 174 510 175
rect 510 174 511 175
rect 511 174 512 175
rect 512 174 513 175
rect 513 174 514 175
rect 514 174 515 175
rect 515 174 516 175
rect 516 174 517 175
rect 517 174 518 175
rect 518 174 519 175
rect 519 174 520 175
rect 102 173 103 174
rect 103 173 104 174
rect 104 173 105 174
rect 105 173 106 174
rect 106 173 107 174
rect 107 173 108 174
rect 108 173 109 174
rect 109 173 110 174
rect 216 173 217 174
rect 217 173 218 174
rect 218 173 219 174
rect 219 173 220 174
rect 220 173 221 174
rect 229 173 230 174
rect 230 173 231 174
rect 231 173 232 174
rect 232 173 233 174
rect 233 173 234 174
rect 234 173 235 174
rect 235 173 236 174
rect 236 173 237 174
rect 237 173 238 174
rect 238 173 239 174
rect 239 173 240 174
rect 240 173 241 174
rect 285 173 286 174
rect 286 173 287 174
rect 287 173 288 174
rect 288 173 289 174
rect 289 173 290 174
rect 290 173 291 174
rect 291 173 292 174
rect 292 173 293 174
rect 293 173 294 174
rect 294 173 295 174
rect 295 173 296 174
rect 296 173 297 174
rect 297 173 298 174
rect 298 173 299 174
rect 330 173 331 174
rect 331 173 332 174
rect 332 173 333 174
rect 333 173 334 174
rect 334 173 335 174
rect 335 173 336 174
rect 336 173 337 174
rect 337 173 338 174
rect 338 173 339 174
rect 339 173 340 174
rect 340 173 341 174
rect 341 173 342 174
rect 342 173 343 174
rect 343 173 344 174
rect 344 173 345 174
rect 345 173 346 174
rect 346 173 347 174
rect 347 173 348 174
rect 348 173 349 174
rect 349 173 350 174
rect 350 173 351 174
rect 351 173 352 174
rect 352 173 353 174
rect 353 173 354 174
rect 375 173 376 174
rect 376 173 377 174
rect 377 173 378 174
rect 378 173 379 174
rect 379 173 380 174
rect 380 173 381 174
rect 381 173 382 174
rect 382 173 383 174
rect 383 173 384 174
rect 384 173 385 174
rect 385 173 386 174
rect 386 173 387 174
rect 387 173 388 174
rect 388 173 389 174
rect 435 173 436 174
rect 436 173 437 174
rect 437 173 438 174
rect 438 173 439 174
rect 439 173 440 174
rect 440 173 441 174
rect 441 173 442 174
rect 442 173 443 174
rect 443 173 444 174
rect 444 173 445 174
rect 504 173 505 174
rect 505 173 506 174
rect 506 173 507 174
rect 507 173 508 174
rect 508 173 509 174
rect 509 173 510 174
rect 510 173 511 174
rect 511 173 512 174
rect 512 173 513 174
rect 513 173 514 174
rect 514 173 515 174
rect 515 173 516 174
rect 516 173 517 174
rect 517 173 518 174
rect 518 173 519 174
rect 519 173 520 174
rect 102 172 103 173
rect 103 172 104 173
rect 104 172 105 173
rect 105 172 106 173
rect 106 172 107 173
rect 107 172 108 173
rect 108 172 109 173
rect 109 172 110 173
rect 110 172 111 173
rect 111 172 112 173
rect 214 172 215 173
rect 215 172 216 173
rect 216 172 217 173
rect 217 172 218 173
rect 218 172 219 173
rect 219 172 220 173
rect 220 172 221 173
rect 229 172 230 173
rect 230 172 231 173
rect 231 172 232 173
rect 232 172 233 173
rect 233 172 234 173
rect 234 172 235 173
rect 235 172 236 173
rect 236 172 237 173
rect 237 172 238 173
rect 238 172 239 173
rect 239 172 240 173
rect 240 172 241 173
rect 283 172 284 173
rect 284 172 285 173
rect 285 172 286 173
rect 286 172 287 173
rect 287 172 288 173
rect 288 172 289 173
rect 289 172 290 173
rect 290 172 291 173
rect 291 172 292 173
rect 292 172 293 173
rect 293 172 294 173
rect 294 172 295 173
rect 295 172 296 173
rect 296 172 297 173
rect 297 172 298 173
rect 298 172 299 173
rect 330 172 331 173
rect 331 172 332 173
rect 332 172 333 173
rect 333 172 334 173
rect 334 172 335 173
rect 335 172 336 173
rect 336 172 337 173
rect 337 172 338 173
rect 338 172 339 173
rect 339 172 340 173
rect 340 172 341 173
rect 341 172 342 173
rect 342 172 343 173
rect 343 172 344 173
rect 344 172 345 173
rect 345 172 346 173
rect 346 172 347 173
rect 347 172 348 173
rect 348 172 349 173
rect 349 172 350 173
rect 350 172 351 173
rect 351 172 352 173
rect 352 172 353 173
rect 353 172 354 173
rect 375 172 376 173
rect 376 172 377 173
rect 377 172 378 173
rect 378 172 379 173
rect 379 172 380 173
rect 380 172 381 173
rect 381 172 382 173
rect 382 172 383 173
rect 383 172 384 173
rect 384 172 385 173
rect 385 172 386 173
rect 386 172 387 173
rect 387 172 388 173
rect 388 172 389 173
rect 389 172 390 173
rect 390 172 391 173
rect 433 172 434 173
rect 434 172 435 173
rect 435 172 436 173
rect 436 172 437 173
rect 437 172 438 173
rect 438 172 439 173
rect 439 172 440 173
rect 440 172 441 173
rect 441 172 442 173
rect 442 172 443 173
rect 443 172 444 173
rect 444 172 445 173
rect 445 172 446 173
rect 446 172 447 173
rect 502 172 503 173
rect 503 172 504 173
rect 504 172 505 173
rect 505 172 506 173
rect 506 172 507 173
rect 507 172 508 173
rect 508 172 509 173
rect 509 172 510 173
rect 510 172 511 173
rect 511 172 512 173
rect 512 172 513 173
rect 513 172 514 173
rect 514 172 515 173
rect 515 172 516 173
rect 516 172 517 173
rect 517 172 518 173
rect 518 172 519 173
rect 519 172 520 173
rect 102 171 103 172
rect 103 171 104 172
rect 104 171 105 172
rect 105 171 106 172
rect 106 171 107 172
rect 107 171 108 172
rect 108 171 109 172
rect 109 171 110 172
rect 110 171 111 172
rect 111 171 112 172
rect 214 171 215 172
rect 215 171 216 172
rect 216 171 217 172
rect 217 171 218 172
rect 218 171 219 172
rect 219 171 220 172
rect 220 171 221 172
rect 231 171 232 172
rect 232 171 233 172
rect 233 171 234 172
rect 234 171 235 172
rect 235 171 236 172
rect 236 171 237 172
rect 237 171 238 172
rect 238 171 239 172
rect 239 171 240 172
rect 240 171 241 172
rect 283 171 284 172
rect 284 171 285 172
rect 285 171 286 172
rect 286 171 287 172
rect 287 171 288 172
rect 288 171 289 172
rect 289 171 290 172
rect 290 171 291 172
rect 291 171 292 172
rect 292 171 293 172
rect 293 171 294 172
rect 294 171 295 172
rect 295 171 296 172
rect 296 171 297 172
rect 297 171 298 172
rect 298 171 299 172
rect 336 171 337 172
rect 337 171 338 172
rect 338 171 339 172
rect 339 171 340 172
rect 340 171 341 172
rect 341 171 342 172
rect 342 171 343 172
rect 343 171 344 172
rect 344 171 345 172
rect 345 171 346 172
rect 346 171 347 172
rect 347 171 348 172
rect 377 171 378 172
rect 378 171 379 172
rect 379 171 380 172
rect 380 171 381 172
rect 381 171 382 172
rect 382 171 383 172
rect 383 171 384 172
rect 384 171 385 172
rect 385 171 386 172
rect 386 171 387 172
rect 387 171 388 172
rect 388 171 389 172
rect 389 171 390 172
rect 390 171 391 172
rect 433 171 434 172
rect 434 171 435 172
rect 435 171 436 172
rect 436 171 437 172
rect 437 171 438 172
rect 438 171 439 172
rect 439 171 440 172
rect 440 171 441 172
rect 441 171 442 172
rect 442 171 443 172
rect 443 171 444 172
rect 444 171 445 172
rect 445 171 446 172
rect 446 171 447 172
rect 502 171 503 172
rect 503 171 504 172
rect 504 171 505 172
rect 505 171 506 172
rect 506 171 507 172
rect 507 171 508 172
rect 508 171 509 172
rect 509 171 510 172
rect 510 171 511 172
rect 511 171 512 172
rect 512 171 513 172
rect 513 171 514 172
rect 514 171 515 172
rect 515 171 516 172
rect 516 171 517 172
rect 517 171 518 172
rect 518 171 519 172
rect 519 171 520 172
rect 102 170 103 171
rect 103 170 104 171
rect 104 170 105 171
rect 105 170 106 171
rect 106 170 107 171
rect 107 170 108 171
rect 108 170 109 171
rect 109 170 110 171
rect 110 170 111 171
rect 111 170 112 171
rect 214 170 215 171
rect 215 170 216 171
rect 216 170 217 171
rect 217 170 218 171
rect 218 170 219 171
rect 219 170 220 171
rect 220 170 221 171
rect 231 170 232 171
rect 232 170 233 171
rect 233 170 234 171
rect 234 170 235 171
rect 235 170 236 171
rect 236 170 237 171
rect 237 170 238 171
rect 238 170 239 171
rect 239 170 240 171
rect 240 170 241 171
rect 241 170 242 171
rect 242 170 243 171
rect 283 170 284 171
rect 284 170 285 171
rect 285 170 286 171
rect 286 170 287 171
rect 287 170 288 171
rect 288 170 289 171
rect 289 170 290 171
rect 290 170 291 171
rect 291 170 292 171
rect 292 170 293 171
rect 293 170 294 171
rect 294 170 295 171
rect 295 170 296 171
rect 296 170 297 171
rect 297 170 298 171
rect 298 170 299 171
rect 299 170 300 171
rect 300 170 301 171
rect 336 170 337 171
rect 337 170 338 171
rect 338 170 339 171
rect 339 170 340 171
rect 340 170 341 171
rect 341 170 342 171
rect 342 170 343 171
rect 343 170 344 171
rect 344 170 345 171
rect 345 170 346 171
rect 346 170 347 171
rect 347 170 348 171
rect 377 170 378 171
rect 378 170 379 171
rect 379 170 380 171
rect 380 170 381 171
rect 381 170 382 171
rect 382 170 383 171
rect 383 170 384 171
rect 384 170 385 171
rect 385 170 386 171
rect 386 170 387 171
rect 387 170 388 171
rect 388 170 389 171
rect 389 170 390 171
rect 390 170 391 171
rect 431 170 432 171
rect 432 170 433 171
rect 433 170 434 171
rect 434 170 435 171
rect 435 170 436 171
rect 436 170 437 171
rect 437 170 438 171
rect 438 170 439 171
rect 439 170 440 171
rect 440 170 441 171
rect 441 170 442 171
rect 442 170 443 171
rect 443 170 444 171
rect 444 170 445 171
rect 445 170 446 171
rect 446 170 447 171
rect 447 170 448 171
rect 448 170 449 171
rect 501 170 502 171
rect 502 170 503 171
rect 503 170 504 171
rect 504 170 505 171
rect 505 170 506 171
rect 506 170 507 171
rect 507 170 508 171
rect 508 170 509 171
rect 509 170 510 171
rect 510 170 511 171
rect 511 170 512 171
rect 512 170 513 171
rect 513 170 514 171
rect 514 170 515 171
rect 515 170 516 171
rect 516 170 517 171
rect 517 170 518 171
rect 518 170 519 171
rect 519 170 520 171
rect 102 169 103 170
rect 103 169 104 170
rect 104 169 105 170
rect 105 169 106 170
rect 106 169 107 170
rect 107 169 108 170
rect 108 169 109 170
rect 109 169 110 170
rect 110 169 111 170
rect 111 169 112 170
rect 214 169 215 170
rect 215 169 216 170
rect 216 169 217 170
rect 217 169 218 170
rect 218 169 219 170
rect 219 169 220 170
rect 220 169 221 170
rect 231 169 232 170
rect 232 169 233 170
rect 233 169 234 170
rect 234 169 235 170
rect 235 169 236 170
rect 236 169 237 170
rect 237 169 238 170
rect 238 169 239 170
rect 239 169 240 170
rect 240 169 241 170
rect 241 169 242 170
rect 242 169 243 170
rect 283 169 284 170
rect 284 169 285 170
rect 285 169 286 170
rect 286 169 287 170
rect 287 169 288 170
rect 289 169 290 170
rect 290 169 291 170
rect 291 169 292 170
rect 292 169 293 170
rect 293 169 294 170
rect 294 169 295 170
rect 295 169 296 170
rect 296 169 297 170
rect 297 169 298 170
rect 298 169 299 170
rect 299 169 300 170
rect 300 169 301 170
rect 336 169 337 170
rect 337 169 338 170
rect 338 169 339 170
rect 339 169 340 170
rect 340 169 341 170
rect 341 169 342 170
rect 342 169 343 170
rect 343 169 344 170
rect 344 169 345 170
rect 345 169 346 170
rect 346 169 347 170
rect 347 169 348 170
rect 379 169 380 170
rect 380 169 381 170
rect 381 169 382 170
rect 382 169 383 170
rect 383 169 384 170
rect 384 169 385 170
rect 385 169 386 170
rect 386 169 387 170
rect 387 169 388 170
rect 388 169 389 170
rect 389 169 390 170
rect 390 169 391 170
rect 431 169 432 170
rect 432 169 433 170
rect 433 169 434 170
rect 434 169 435 170
rect 435 169 436 170
rect 436 169 437 170
rect 437 169 438 170
rect 438 169 439 170
rect 439 169 440 170
rect 440 169 441 170
rect 441 169 442 170
rect 442 169 443 170
rect 443 169 444 170
rect 444 169 445 170
rect 445 169 446 170
rect 446 169 447 170
rect 447 169 448 170
rect 448 169 449 170
rect 501 169 502 170
rect 502 169 503 170
rect 503 169 504 170
rect 504 169 505 170
rect 505 169 506 170
rect 506 169 507 170
rect 507 169 508 170
rect 508 169 509 170
rect 509 169 510 170
rect 510 169 511 170
rect 511 169 512 170
rect 512 169 513 170
rect 513 169 514 170
rect 514 169 515 170
rect 515 169 516 170
rect 516 169 517 170
rect 517 169 518 170
rect 102 168 103 169
rect 103 168 104 169
rect 104 168 105 169
rect 105 168 106 169
rect 106 168 107 169
rect 107 168 108 169
rect 108 168 109 169
rect 109 168 110 169
rect 110 168 111 169
rect 111 168 112 169
rect 112 168 113 169
rect 113 168 114 169
rect 214 168 215 169
rect 215 168 216 169
rect 216 168 217 169
rect 217 168 218 169
rect 218 168 219 169
rect 219 168 220 169
rect 220 168 221 169
rect 231 168 232 169
rect 232 168 233 169
rect 233 168 234 169
rect 234 168 235 169
rect 235 168 236 169
rect 236 168 237 169
rect 237 168 238 169
rect 238 168 239 169
rect 239 168 240 169
rect 240 168 241 169
rect 241 168 242 169
rect 242 168 243 169
rect 281 168 282 169
rect 282 168 283 169
rect 283 168 284 169
rect 284 168 285 169
rect 285 168 286 169
rect 286 168 287 169
rect 287 168 288 169
rect 289 168 290 169
rect 290 168 291 169
rect 291 168 292 169
rect 292 168 293 169
rect 293 168 294 169
rect 294 168 295 169
rect 295 168 296 169
rect 296 168 297 169
rect 297 168 298 169
rect 298 168 299 169
rect 299 168 300 169
rect 300 168 301 169
rect 336 168 337 169
rect 337 168 338 169
rect 338 168 339 169
rect 339 168 340 169
rect 340 168 341 169
rect 341 168 342 169
rect 342 168 343 169
rect 343 168 344 169
rect 344 168 345 169
rect 345 168 346 169
rect 346 168 347 169
rect 347 168 348 169
rect 379 168 380 169
rect 380 168 381 169
rect 381 168 382 169
rect 382 168 383 169
rect 383 168 384 169
rect 384 168 385 169
rect 385 168 386 169
rect 386 168 387 169
rect 387 168 388 169
rect 388 168 389 169
rect 389 168 390 169
rect 390 168 391 169
rect 391 168 392 169
rect 392 168 393 169
rect 426 168 427 169
rect 427 168 428 169
rect 428 168 429 169
rect 429 168 430 169
rect 430 168 431 169
rect 431 168 432 169
rect 432 168 433 169
rect 433 168 434 169
rect 434 168 435 169
rect 435 168 436 169
rect 436 168 437 169
rect 437 168 438 169
rect 438 168 439 169
rect 439 168 440 169
rect 440 168 441 169
rect 441 168 442 169
rect 442 168 443 169
rect 443 168 444 169
rect 444 168 445 169
rect 445 168 446 169
rect 446 168 447 169
rect 447 168 448 169
rect 448 168 449 169
rect 449 168 450 169
rect 450 168 451 169
rect 451 168 452 169
rect 452 168 453 169
rect 453 168 454 169
rect 454 168 455 169
rect 501 168 502 169
rect 502 168 503 169
rect 503 168 504 169
rect 504 168 505 169
rect 505 168 506 169
rect 506 168 507 169
rect 507 168 508 169
rect 508 168 509 169
rect 509 168 510 169
rect 510 168 511 169
rect 511 168 512 169
rect 512 168 513 169
rect 513 168 514 169
rect 514 168 515 169
rect 515 168 516 169
rect 516 168 517 169
rect 517 168 518 169
rect 103 167 104 168
rect 104 167 105 168
rect 105 167 106 168
rect 106 167 107 168
rect 107 167 108 168
rect 108 167 109 168
rect 109 167 110 168
rect 110 167 111 168
rect 111 167 112 168
rect 112 167 113 168
rect 113 167 114 168
rect 214 167 215 168
rect 215 167 216 168
rect 216 167 217 168
rect 217 167 218 168
rect 218 167 219 168
rect 231 167 232 168
rect 232 167 233 168
rect 233 167 234 168
rect 234 167 235 168
rect 235 167 236 168
rect 236 167 237 168
rect 237 167 238 168
rect 238 167 239 168
rect 239 167 240 168
rect 240 167 241 168
rect 241 167 242 168
rect 242 167 243 168
rect 281 167 282 168
rect 282 167 283 168
rect 283 167 284 168
rect 284 167 285 168
rect 285 167 286 168
rect 286 167 287 168
rect 287 167 288 168
rect 289 167 290 168
rect 290 167 291 168
rect 291 167 292 168
rect 292 167 293 168
rect 293 167 294 168
rect 294 167 295 168
rect 295 167 296 168
rect 296 167 297 168
rect 297 167 298 168
rect 298 167 299 168
rect 299 167 300 168
rect 300 167 301 168
rect 336 167 337 168
rect 337 167 338 168
rect 338 167 339 168
rect 339 167 340 168
rect 340 167 341 168
rect 341 167 342 168
rect 342 167 343 168
rect 343 167 344 168
rect 344 167 345 168
rect 345 167 346 168
rect 379 167 380 168
rect 380 167 381 168
rect 381 167 382 168
rect 382 167 383 168
rect 383 167 384 168
rect 384 167 385 168
rect 385 167 386 168
rect 386 167 387 168
rect 387 167 388 168
rect 388 167 389 168
rect 389 167 390 168
rect 390 167 391 168
rect 391 167 392 168
rect 392 167 393 168
rect 426 167 427 168
rect 427 167 428 168
rect 428 167 429 168
rect 429 167 430 168
rect 430 167 431 168
rect 431 167 432 168
rect 432 167 433 168
rect 433 167 434 168
rect 434 167 435 168
rect 435 167 436 168
rect 436 167 437 168
rect 437 167 438 168
rect 438 167 439 168
rect 439 167 440 168
rect 440 167 441 168
rect 441 167 442 168
rect 442 167 443 168
rect 443 167 444 168
rect 444 167 445 168
rect 445 167 446 168
rect 446 167 447 168
rect 447 167 448 168
rect 448 167 449 168
rect 449 167 450 168
rect 450 167 451 168
rect 451 167 452 168
rect 452 167 453 168
rect 453 167 454 168
rect 454 167 455 168
rect 501 167 502 168
rect 502 167 503 168
rect 503 167 504 168
rect 504 167 505 168
rect 505 167 506 168
rect 506 167 507 168
rect 507 167 508 168
rect 508 167 509 168
rect 509 167 510 168
rect 510 167 511 168
rect 511 167 512 168
rect 512 167 513 168
rect 513 167 514 168
rect 514 167 515 168
rect 515 167 516 168
rect 516 167 517 168
rect 517 167 518 168
rect 103 166 104 167
rect 104 166 105 167
rect 105 166 106 167
rect 106 166 107 167
rect 107 166 108 167
rect 108 166 109 167
rect 109 166 110 167
rect 110 166 111 167
rect 111 166 112 167
rect 112 166 113 167
rect 113 166 114 167
rect 212 166 213 167
rect 213 166 214 167
rect 214 166 215 167
rect 215 166 216 167
rect 216 166 217 167
rect 217 166 218 167
rect 218 166 219 167
rect 231 166 232 167
rect 232 166 233 167
rect 233 166 234 167
rect 234 166 235 167
rect 235 166 236 167
rect 236 166 237 167
rect 237 166 238 167
rect 238 166 239 167
rect 239 166 240 167
rect 240 166 241 167
rect 241 166 242 167
rect 242 166 243 167
rect 243 166 244 167
rect 244 166 245 167
rect 281 166 282 167
rect 282 166 283 167
rect 283 166 284 167
rect 284 166 285 167
rect 285 166 286 167
rect 286 166 287 167
rect 287 166 288 167
rect 289 166 290 167
rect 290 166 291 167
rect 291 166 292 167
rect 292 166 293 167
rect 293 166 294 167
rect 294 166 295 167
rect 295 166 296 167
rect 296 166 297 167
rect 297 166 298 167
rect 298 166 299 167
rect 299 166 300 167
rect 300 166 301 167
rect 336 166 337 167
rect 337 166 338 167
rect 338 166 339 167
rect 339 166 340 167
rect 340 166 341 167
rect 341 166 342 167
rect 342 166 343 167
rect 343 166 344 167
rect 344 166 345 167
rect 345 166 346 167
rect 379 166 380 167
rect 380 166 381 167
rect 381 166 382 167
rect 382 166 383 167
rect 383 166 384 167
rect 384 166 385 167
rect 385 166 386 167
rect 386 166 387 167
rect 387 166 388 167
rect 388 166 389 167
rect 389 166 390 167
rect 390 166 391 167
rect 391 166 392 167
rect 392 166 393 167
rect 426 166 427 167
rect 427 166 428 167
rect 428 166 429 167
rect 429 166 430 167
rect 430 166 431 167
rect 431 166 432 167
rect 432 166 433 167
rect 433 166 434 167
rect 434 166 435 167
rect 435 166 436 167
rect 436 166 437 167
rect 437 166 438 167
rect 438 166 439 167
rect 439 166 440 167
rect 440 166 441 167
rect 441 166 442 167
rect 442 166 443 167
rect 443 166 444 167
rect 444 166 445 167
rect 445 166 446 167
rect 446 166 447 167
rect 447 166 448 167
rect 448 166 449 167
rect 449 166 450 167
rect 450 166 451 167
rect 451 166 452 167
rect 452 166 453 167
rect 453 166 454 167
rect 454 166 455 167
rect 499 166 500 167
rect 500 166 501 167
rect 501 166 502 167
rect 502 166 503 167
rect 503 166 504 167
rect 504 166 505 167
rect 505 166 506 167
rect 506 166 507 167
rect 507 166 508 167
rect 508 166 509 167
rect 509 166 510 167
rect 510 166 511 167
rect 511 166 512 167
rect 512 166 513 167
rect 513 166 514 167
rect 514 166 515 167
rect 515 166 516 167
rect 516 166 517 167
rect 517 166 518 167
rect 103 165 104 166
rect 104 165 105 166
rect 105 165 106 166
rect 106 165 107 166
rect 107 165 108 166
rect 108 165 109 166
rect 109 165 110 166
rect 110 165 111 166
rect 111 165 112 166
rect 112 165 113 166
rect 113 165 114 166
rect 212 165 213 166
rect 213 165 214 166
rect 214 165 215 166
rect 215 165 216 166
rect 216 165 217 166
rect 217 165 218 166
rect 218 165 219 166
rect 233 165 234 166
rect 234 165 235 166
rect 235 165 236 166
rect 236 165 237 166
rect 237 165 238 166
rect 238 165 239 166
rect 239 165 240 166
rect 240 165 241 166
rect 241 165 242 166
rect 242 165 243 166
rect 243 165 244 166
rect 244 165 245 166
rect 281 165 282 166
rect 282 165 283 166
rect 283 165 284 166
rect 284 165 285 166
rect 285 165 286 166
rect 286 165 287 166
rect 287 165 288 166
rect 291 165 292 166
rect 292 165 293 166
rect 293 165 294 166
rect 294 165 295 166
rect 295 165 296 166
rect 296 165 297 166
rect 297 165 298 166
rect 298 165 299 166
rect 299 165 300 166
rect 300 165 301 166
rect 336 165 337 166
rect 337 165 338 166
rect 338 165 339 166
rect 339 165 340 166
rect 340 165 341 166
rect 341 165 342 166
rect 342 165 343 166
rect 343 165 344 166
rect 344 165 345 166
rect 345 165 346 166
rect 381 165 382 166
rect 382 165 383 166
rect 383 165 384 166
rect 384 165 385 166
rect 385 165 386 166
rect 386 165 387 166
rect 387 165 388 166
rect 388 165 389 166
rect 389 165 390 166
rect 390 165 391 166
rect 391 165 392 166
rect 392 165 393 166
rect 499 165 500 166
rect 500 165 501 166
rect 501 165 502 166
rect 502 165 503 166
rect 503 165 504 166
rect 504 165 505 166
rect 505 165 506 166
rect 506 165 507 166
rect 507 165 508 166
rect 508 165 509 166
rect 509 165 510 166
rect 510 165 511 166
rect 511 165 512 166
rect 512 165 513 166
rect 513 165 514 166
rect 514 165 515 166
rect 515 165 516 166
rect 103 164 104 165
rect 104 164 105 165
rect 105 164 106 165
rect 106 164 107 165
rect 107 164 108 165
rect 108 164 109 165
rect 109 164 110 165
rect 110 164 111 165
rect 111 164 112 165
rect 112 164 113 165
rect 113 164 114 165
rect 114 164 115 165
rect 115 164 116 165
rect 212 164 213 165
rect 213 164 214 165
rect 214 164 215 165
rect 215 164 216 165
rect 216 164 217 165
rect 217 164 218 165
rect 218 164 219 165
rect 233 164 234 165
rect 234 164 235 165
rect 235 164 236 165
rect 236 164 237 165
rect 237 164 238 165
rect 238 164 239 165
rect 239 164 240 165
rect 240 164 241 165
rect 241 164 242 165
rect 242 164 243 165
rect 243 164 244 165
rect 244 164 245 165
rect 281 164 282 165
rect 282 164 283 165
rect 283 164 284 165
rect 284 164 285 165
rect 285 164 286 165
rect 286 164 287 165
rect 287 164 288 165
rect 291 164 292 165
rect 292 164 293 165
rect 293 164 294 165
rect 294 164 295 165
rect 295 164 296 165
rect 296 164 297 165
rect 297 164 298 165
rect 298 164 299 165
rect 299 164 300 165
rect 300 164 301 165
rect 301 164 302 165
rect 302 164 303 165
rect 336 164 337 165
rect 337 164 338 165
rect 338 164 339 165
rect 339 164 340 165
rect 340 164 341 165
rect 341 164 342 165
rect 342 164 343 165
rect 343 164 344 165
rect 344 164 345 165
rect 345 164 346 165
rect 346 164 347 165
rect 347 164 348 165
rect 381 164 382 165
rect 382 164 383 165
rect 383 164 384 165
rect 384 164 385 165
rect 385 164 386 165
rect 386 164 387 165
rect 387 164 388 165
rect 388 164 389 165
rect 389 164 390 165
rect 390 164 391 165
rect 391 164 392 165
rect 392 164 393 165
rect 497 164 498 165
rect 498 164 499 165
rect 499 164 500 165
rect 500 164 501 165
rect 501 164 502 165
rect 502 164 503 165
rect 503 164 504 165
rect 504 164 505 165
rect 505 164 506 165
rect 506 164 507 165
rect 507 164 508 165
rect 508 164 509 165
rect 509 164 510 165
rect 510 164 511 165
rect 511 164 512 165
rect 512 164 513 165
rect 513 164 514 165
rect 514 164 515 165
rect 515 164 516 165
rect 105 163 106 164
rect 106 163 107 164
rect 107 163 108 164
rect 108 163 109 164
rect 109 163 110 164
rect 110 163 111 164
rect 111 163 112 164
rect 112 163 113 164
rect 113 163 114 164
rect 114 163 115 164
rect 115 163 116 164
rect 212 163 213 164
rect 213 163 214 164
rect 214 163 215 164
rect 215 163 216 164
rect 216 163 217 164
rect 217 163 218 164
rect 218 163 219 164
rect 233 163 234 164
rect 234 163 235 164
rect 235 163 236 164
rect 236 163 237 164
rect 237 163 238 164
rect 238 163 239 164
rect 239 163 240 164
rect 240 163 241 164
rect 241 163 242 164
rect 242 163 243 164
rect 243 163 244 164
rect 244 163 245 164
rect 281 163 282 164
rect 282 163 283 164
rect 283 163 284 164
rect 284 163 285 164
rect 285 163 286 164
rect 291 163 292 164
rect 292 163 293 164
rect 293 163 294 164
rect 294 163 295 164
rect 295 163 296 164
rect 296 163 297 164
rect 297 163 298 164
rect 298 163 299 164
rect 299 163 300 164
rect 300 163 301 164
rect 301 163 302 164
rect 302 163 303 164
rect 336 163 337 164
rect 337 163 338 164
rect 338 163 339 164
rect 339 163 340 164
rect 340 163 341 164
rect 341 163 342 164
rect 342 163 343 164
rect 343 163 344 164
rect 344 163 345 164
rect 345 163 346 164
rect 346 163 347 164
rect 347 163 348 164
rect 383 163 384 164
rect 384 163 385 164
rect 385 163 386 164
rect 386 163 387 164
rect 387 163 388 164
rect 388 163 389 164
rect 389 163 390 164
rect 390 163 391 164
rect 497 163 498 164
rect 498 163 499 164
rect 499 163 500 164
rect 500 163 501 164
rect 501 163 502 164
rect 502 163 503 164
rect 503 163 504 164
rect 504 163 505 164
rect 505 163 506 164
rect 506 163 507 164
rect 507 163 508 164
rect 508 163 509 164
rect 509 163 510 164
rect 510 163 511 164
rect 511 163 512 164
rect 512 163 513 164
rect 513 163 514 164
rect 514 163 515 164
rect 515 163 516 164
rect 105 162 106 163
rect 106 162 107 163
rect 107 162 108 163
rect 108 162 109 163
rect 109 162 110 163
rect 110 162 111 163
rect 111 162 112 163
rect 112 162 113 163
rect 113 162 114 163
rect 114 162 115 163
rect 115 162 116 163
rect 212 162 213 163
rect 213 162 214 163
rect 214 162 215 163
rect 215 162 216 163
rect 216 162 217 163
rect 217 162 218 163
rect 218 162 219 163
rect 233 162 234 163
rect 234 162 235 163
rect 235 162 236 163
rect 236 162 237 163
rect 237 162 238 163
rect 238 162 239 163
rect 239 162 240 163
rect 240 162 241 163
rect 241 162 242 163
rect 242 162 243 163
rect 243 162 244 163
rect 244 162 245 163
rect 279 162 280 163
rect 280 162 281 163
rect 281 162 282 163
rect 282 162 283 163
rect 283 162 284 163
rect 284 162 285 163
rect 285 162 286 163
rect 291 162 292 163
rect 292 162 293 163
rect 293 162 294 163
rect 294 162 295 163
rect 295 162 296 163
rect 296 162 297 163
rect 297 162 298 163
rect 298 162 299 163
rect 299 162 300 163
rect 300 162 301 163
rect 301 162 302 163
rect 302 162 303 163
rect 336 162 337 163
rect 337 162 338 163
rect 338 162 339 163
rect 339 162 340 163
rect 340 162 341 163
rect 341 162 342 163
rect 342 162 343 163
rect 343 162 344 163
rect 344 162 345 163
rect 345 162 346 163
rect 346 162 347 163
rect 347 162 348 163
rect 383 162 384 163
rect 384 162 385 163
rect 385 162 386 163
rect 386 162 387 163
rect 387 162 388 163
rect 388 162 389 163
rect 389 162 390 163
rect 390 162 391 163
rect 495 162 496 163
rect 496 162 497 163
rect 497 162 498 163
rect 498 162 499 163
rect 499 162 500 163
rect 500 162 501 163
rect 501 162 502 163
rect 502 162 503 163
rect 503 162 504 163
rect 504 162 505 163
rect 505 162 506 163
rect 506 162 507 163
rect 507 162 508 163
rect 508 162 509 163
rect 509 162 510 163
rect 510 162 511 163
rect 511 162 512 163
rect 512 162 513 163
rect 513 162 514 163
rect 514 162 515 163
rect 515 162 516 163
rect 105 161 106 162
rect 106 161 107 162
rect 107 161 108 162
rect 108 161 109 162
rect 109 161 110 162
rect 110 161 111 162
rect 111 161 112 162
rect 112 161 113 162
rect 113 161 114 162
rect 114 161 115 162
rect 115 161 116 162
rect 212 161 213 162
rect 213 161 214 162
rect 214 161 215 162
rect 215 161 216 162
rect 216 161 217 162
rect 235 161 236 162
rect 236 161 237 162
rect 237 161 238 162
rect 238 161 239 162
rect 239 161 240 162
rect 240 161 241 162
rect 241 161 242 162
rect 242 161 243 162
rect 243 161 244 162
rect 244 161 245 162
rect 279 161 280 162
rect 280 161 281 162
rect 281 161 282 162
rect 282 161 283 162
rect 283 161 284 162
rect 284 161 285 162
rect 285 161 286 162
rect 293 161 294 162
rect 294 161 295 162
rect 295 161 296 162
rect 296 161 297 162
rect 297 161 298 162
rect 298 161 299 162
rect 299 161 300 162
rect 300 161 301 162
rect 301 161 302 162
rect 302 161 303 162
rect 336 161 337 162
rect 337 161 338 162
rect 338 161 339 162
rect 339 161 340 162
rect 340 161 341 162
rect 341 161 342 162
rect 342 161 343 162
rect 343 161 344 162
rect 344 161 345 162
rect 345 161 346 162
rect 383 161 384 162
rect 384 161 385 162
rect 385 161 386 162
rect 386 161 387 162
rect 387 161 388 162
rect 388 161 389 162
rect 495 161 496 162
rect 496 161 497 162
rect 497 161 498 162
rect 498 161 499 162
rect 499 161 500 162
rect 500 161 501 162
rect 501 161 502 162
rect 502 161 503 162
rect 503 161 504 162
rect 504 161 505 162
rect 505 161 506 162
rect 506 161 507 162
rect 507 161 508 162
rect 508 161 509 162
rect 509 161 510 162
rect 510 161 511 162
rect 511 161 512 162
rect 512 161 513 162
rect 513 161 514 162
rect 514 161 515 162
rect 105 160 106 161
rect 106 160 107 161
rect 107 160 108 161
rect 108 160 109 161
rect 109 160 110 161
rect 110 160 111 161
rect 111 160 112 161
rect 112 160 113 161
rect 113 160 114 161
rect 114 160 115 161
rect 115 160 116 161
rect 116 160 117 161
rect 117 160 118 161
rect 210 160 211 161
rect 211 160 212 161
rect 212 160 213 161
rect 213 160 214 161
rect 214 160 215 161
rect 215 160 216 161
rect 216 160 217 161
rect 235 160 236 161
rect 236 160 237 161
rect 237 160 238 161
rect 238 160 239 161
rect 239 160 240 161
rect 240 160 241 161
rect 241 160 242 161
rect 242 160 243 161
rect 243 160 244 161
rect 244 160 245 161
rect 245 160 246 161
rect 246 160 247 161
rect 279 160 280 161
rect 280 160 281 161
rect 281 160 282 161
rect 282 160 283 161
rect 283 160 284 161
rect 284 160 285 161
rect 285 160 286 161
rect 293 160 294 161
rect 294 160 295 161
rect 295 160 296 161
rect 296 160 297 161
rect 297 160 298 161
rect 298 160 299 161
rect 299 160 300 161
rect 300 160 301 161
rect 301 160 302 161
rect 302 160 303 161
rect 303 160 304 161
rect 304 160 305 161
rect 336 160 337 161
rect 337 160 338 161
rect 338 160 339 161
rect 339 160 340 161
rect 340 160 341 161
rect 341 160 342 161
rect 342 160 343 161
rect 343 160 344 161
rect 344 160 345 161
rect 345 160 346 161
rect 381 160 382 161
rect 382 160 383 161
rect 383 160 384 161
rect 384 160 385 161
rect 385 160 386 161
rect 386 160 387 161
rect 387 160 388 161
rect 388 160 389 161
rect 495 160 496 161
rect 496 160 497 161
rect 497 160 498 161
rect 498 160 499 161
rect 499 160 500 161
rect 500 160 501 161
rect 501 160 502 161
rect 502 160 503 161
rect 503 160 504 161
rect 504 160 505 161
rect 505 160 506 161
rect 506 160 507 161
rect 507 160 508 161
rect 508 160 509 161
rect 509 160 510 161
rect 510 160 511 161
rect 511 160 512 161
rect 512 160 513 161
rect 513 160 514 161
rect 514 160 515 161
rect 107 159 108 160
rect 108 159 109 160
rect 109 159 110 160
rect 110 159 111 160
rect 111 159 112 160
rect 112 159 113 160
rect 113 159 114 160
rect 114 159 115 160
rect 115 159 116 160
rect 116 159 117 160
rect 117 159 118 160
rect 210 159 211 160
rect 211 159 212 160
rect 212 159 213 160
rect 213 159 214 160
rect 214 159 215 160
rect 215 159 216 160
rect 216 159 217 160
rect 235 159 236 160
rect 236 159 237 160
rect 237 159 238 160
rect 238 159 239 160
rect 239 159 240 160
rect 240 159 241 160
rect 241 159 242 160
rect 242 159 243 160
rect 243 159 244 160
rect 244 159 245 160
rect 245 159 246 160
rect 246 159 247 160
rect 279 159 280 160
rect 280 159 281 160
rect 281 159 282 160
rect 282 159 283 160
rect 283 159 284 160
rect 284 159 285 160
rect 285 159 286 160
rect 293 159 294 160
rect 294 159 295 160
rect 295 159 296 160
rect 296 159 297 160
rect 297 159 298 160
rect 298 159 299 160
rect 299 159 300 160
rect 300 159 301 160
rect 301 159 302 160
rect 302 159 303 160
rect 303 159 304 160
rect 304 159 305 160
rect 336 159 337 160
rect 337 159 338 160
rect 338 159 339 160
rect 339 159 340 160
rect 340 159 341 160
rect 341 159 342 160
rect 342 159 343 160
rect 343 159 344 160
rect 344 159 345 160
rect 345 159 346 160
rect 381 159 382 160
rect 382 159 383 160
rect 383 159 384 160
rect 384 159 385 160
rect 385 159 386 160
rect 386 159 387 160
rect 387 159 388 160
rect 388 159 389 160
rect 495 159 496 160
rect 496 159 497 160
rect 497 159 498 160
rect 498 159 499 160
rect 499 159 500 160
rect 500 159 501 160
rect 501 159 502 160
rect 502 159 503 160
rect 503 159 504 160
rect 504 159 505 160
rect 505 159 506 160
rect 506 159 507 160
rect 507 159 508 160
rect 508 159 509 160
rect 509 159 510 160
rect 510 159 511 160
rect 511 159 512 160
rect 512 159 513 160
rect 513 159 514 160
rect 514 159 515 160
rect 107 158 108 159
rect 108 158 109 159
rect 109 158 110 159
rect 110 158 111 159
rect 111 158 112 159
rect 112 158 113 159
rect 113 158 114 159
rect 114 158 115 159
rect 115 158 116 159
rect 116 158 117 159
rect 117 158 118 159
rect 210 158 211 159
rect 211 158 212 159
rect 212 158 213 159
rect 213 158 214 159
rect 214 158 215 159
rect 215 158 216 159
rect 216 158 217 159
rect 235 158 236 159
rect 236 158 237 159
rect 237 158 238 159
rect 238 158 239 159
rect 239 158 240 159
rect 240 158 241 159
rect 241 158 242 159
rect 242 158 243 159
rect 243 158 244 159
rect 244 158 245 159
rect 245 158 246 159
rect 246 158 247 159
rect 279 158 280 159
rect 280 158 281 159
rect 281 158 282 159
rect 282 158 283 159
rect 283 158 284 159
rect 284 158 285 159
rect 285 158 286 159
rect 293 158 294 159
rect 294 158 295 159
rect 295 158 296 159
rect 296 158 297 159
rect 297 158 298 159
rect 298 158 299 159
rect 299 158 300 159
rect 300 158 301 159
rect 301 158 302 159
rect 302 158 303 159
rect 303 158 304 159
rect 304 158 305 159
rect 336 158 337 159
rect 337 158 338 159
rect 338 158 339 159
rect 339 158 340 159
rect 340 158 341 159
rect 341 158 342 159
rect 342 158 343 159
rect 343 158 344 159
rect 344 158 345 159
rect 345 158 346 159
rect 381 158 382 159
rect 382 158 383 159
rect 383 158 384 159
rect 384 158 385 159
rect 385 158 386 159
rect 386 158 387 159
rect 387 158 388 159
rect 388 158 389 159
rect 493 158 494 159
rect 494 158 495 159
rect 495 158 496 159
rect 496 158 497 159
rect 497 158 498 159
rect 498 158 499 159
rect 499 158 500 159
rect 500 158 501 159
rect 501 158 502 159
rect 502 158 503 159
rect 503 158 504 159
rect 504 158 505 159
rect 505 158 506 159
rect 506 158 507 159
rect 507 158 508 159
rect 508 158 509 159
rect 509 158 510 159
rect 510 158 511 159
rect 511 158 512 159
rect 512 158 513 159
rect 513 158 514 159
rect 514 158 515 159
rect 107 157 108 158
rect 108 157 109 158
rect 109 157 110 158
rect 110 157 111 158
rect 111 157 112 158
rect 112 157 113 158
rect 113 157 114 158
rect 114 157 115 158
rect 115 157 116 158
rect 116 157 117 158
rect 117 157 118 158
rect 210 157 211 158
rect 211 157 212 158
rect 212 157 213 158
rect 213 157 214 158
rect 214 157 215 158
rect 215 157 216 158
rect 216 157 217 158
rect 235 157 236 158
rect 236 157 237 158
rect 237 157 238 158
rect 238 157 239 158
rect 239 157 240 158
rect 240 157 241 158
rect 241 157 242 158
rect 242 157 243 158
rect 243 157 244 158
rect 244 157 245 158
rect 245 157 246 158
rect 246 157 247 158
rect 279 157 280 158
rect 280 157 281 158
rect 281 157 282 158
rect 282 157 283 158
rect 283 157 284 158
rect 293 157 294 158
rect 294 157 295 158
rect 295 157 296 158
rect 296 157 297 158
rect 297 157 298 158
rect 298 157 299 158
rect 299 157 300 158
rect 300 157 301 158
rect 301 157 302 158
rect 302 157 303 158
rect 303 157 304 158
rect 304 157 305 158
rect 336 157 337 158
rect 337 157 338 158
rect 338 157 339 158
rect 339 157 340 158
rect 340 157 341 158
rect 341 157 342 158
rect 342 157 343 158
rect 343 157 344 158
rect 344 157 345 158
rect 345 157 346 158
rect 381 157 382 158
rect 382 157 383 158
rect 383 157 384 158
rect 384 157 385 158
rect 493 157 494 158
rect 494 157 495 158
rect 495 157 496 158
rect 496 157 497 158
rect 497 157 498 158
rect 498 157 499 158
rect 499 157 500 158
rect 500 157 501 158
rect 501 157 502 158
rect 502 157 503 158
rect 503 157 504 158
rect 504 157 505 158
rect 505 157 506 158
rect 506 157 507 158
rect 507 157 508 158
rect 508 157 509 158
rect 509 157 510 158
rect 510 157 511 158
rect 511 157 512 158
rect 512 157 513 158
rect 107 156 108 157
rect 108 156 109 157
rect 109 156 110 157
rect 110 156 111 157
rect 111 156 112 157
rect 112 156 113 157
rect 113 156 114 157
rect 114 156 115 157
rect 115 156 116 157
rect 116 156 117 157
rect 117 156 118 157
rect 118 156 119 157
rect 208 156 209 157
rect 209 156 210 157
rect 210 156 211 157
rect 211 156 212 157
rect 212 156 213 157
rect 213 156 214 157
rect 214 156 215 157
rect 215 156 216 157
rect 216 156 217 157
rect 235 156 236 157
rect 236 156 237 157
rect 237 156 238 157
rect 238 156 239 157
rect 239 156 240 157
rect 240 156 241 157
rect 241 156 242 157
rect 242 156 243 157
rect 243 156 244 157
rect 244 156 245 157
rect 245 156 246 157
rect 246 156 247 157
rect 247 156 248 157
rect 248 156 249 157
rect 278 156 279 157
rect 279 156 280 157
rect 280 156 281 157
rect 281 156 282 157
rect 282 156 283 157
rect 283 156 284 157
rect 293 156 294 157
rect 294 156 295 157
rect 295 156 296 157
rect 296 156 297 157
rect 297 156 298 157
rect 298 156 299 157
rect 299 156 300 157
rect 300 156 301 157
rect 301 156 302 157
rect 302 156 303 157
rect 303 156 304 157
rect 304 156 305 157
rect 336 156 337 157
rect 337 156 338 157
rect 338 156 339 157
rect 339 156 340 157
rect 340 156 341 157
rect 341 156 342 157
rect 342 156 343 157
rect 343 156 344 157
rect 344 156 345 157
rect 345 156 346 157
rect 346 156 347 157
rect 347 156 348 157
rect 377 156 378 157
rect 378 156 379 157
rect 379 156 380 157
rect 380 156 381 157
rect 381 156 382 157
rect 382 156 383 157
rect 383 156 384 157
rect 384 156 385 157
rect 491 156 492 157
rect 492 156 493 157
rect 493 156 494 157
rect 494 156 495 157
rect 495 156 496 157
rect 496 156 497 157
rect 497 156 498 157
rect 498 156 499 157
rect 499 156 500 157
rect 500 156 501 157
rect 501 156 502 157
rect 502 156 503 157
rect 503 156 504 157
rect 504 156 505 157
rect 505 156 506 157
rect 506 156 507 157
rect 507 156 508 157
rect 508 156 509 157
rect 509 156 510 157
rect 510 156 511 157
rect 511 156 512 157
rect 512 156 513 157
rect 107 155 108 156
rect 108 155 109 156
rect 109 155 110 156
rect 110 155 111 156
rect 111 155 112 156
rect 112 155 113 156
rect 113 155 114 156
rect 114 155 115 156
rect 115 155 116 156
rect 116 155 117 156
rect 117 155 118 156
rect 118 155 119 156
rect 208 155 209 156
rect 209 155 210 156
rect 210 155 211 156
rect 211 155 212 156
rect 212 155 213 156
rect 213 155 214 156
rect 214 155 215 156
rect 236 155 237 156
rect 237 155 238 156
rect 238 155 239 156
rect 239 155 240 156
rect 240 155 241 156
rect 241 155 242 156
rect 242 155 243 156
rect 243 155 244 156
rect 244 155 245 156
rect 245 155 246 156
rect 246 155 247 156
rect 247 155 248 156
rect 248 155 249 156
rect 278 155 279 156
rect 279 155 280 156
rect 280 155 281 156
rect 281 155 282 156
rect 282 155 283 156
rect 283 155 284 156
rect 294 155 295 156
rect 295 155 296 156
rect 296 155 297 156
rect 297 155 298 156
rect 298 155 299 156
rect 299 155 300 156
rect 300 155 301 156
rect 301 155 302 156
rect 302 155 303 156
rect 303 155 304 156
rect 304 155 305 156
rect 336 155 337 156
rect 337 155 338 156
rect 338 155 339 156
rect 339 155 340 156
rect 340 155 341 156
rect 341 155 342 156
rect 342 155 343 156
rect 343 155 344 156
rect 344 155 345 156
rect 345 155 346 156
rect 346 155 347 156
rect 347 155 348 156
rect 377 155 378 156
rect 378 155 379 156
rect 379 155 380 156
rect 380 155 381 156
rect 381 155 382 156
rect 382 155 383 156
rect 383 155 384 156
rect 384 155 385 156
rect 491 155 492 156
rect 492 155 493 156
rect 493 155 494 156
rect 494 155 495 156
rect 495 155 496 156
rect 496 155 497 156
rect 497 155 498 156
rect 498 155 499 156
rect 499 155 500 156
rect 500 155 501 156
rect 501 155 502 156
rect 502 155 503 156
rect 503 155 504 156
rect 504 155 505 156
rect 505 155 506 156
rect 506 155 507 156
rect 507 155 508 156
rect 508 155 509 156
rect 509 155 510 156
rect 510 155 511 156
rect 511 155 512 156
rect 512 155 513 156
rect 107 154 108 155
rect 108 154 109 155
rect 109 154 110 155
rect 110 154 111 155
rect 111 154 112 155
rect 112 154 113 155
rect 113 154 114 155
rect 114 154 115 155
rect 115 154 116 155
rect 116 154 117 155
rect 117 154 118 155
rect 118 154 119 155
rect 208 154 209 155
rect 209 154 210 155
rect 210 154 211 155
rect 211 154 212 155
rect 212 154 213 155
rect 213 154 214 155
rect 214 154 215 155
rect 236 154 237 155
rect 237 154 238 155
rect 238 154 239 155
rect 239 154 240 155
rect 240 154 241 155
rect 241 154 242 155
rect 242 154 243 155
rect 243 154 244 155
rect 244 154 245 155
rect 245 154 246 155
rect 246 154 247 155
rect 247 154 248 155
rect 248 154 249 155
rect 278 154 279 155
rect 279 154 280 155
rect 280 154 281 155
rect 281 154 282 155
rect 282 154 283 155
rect 283 154 284 155
rect 294 154 295 155
rect 295 154 296 155
rect 296 154 297 155
rect 297 154 298 155
rect 298 154 299 155
rect 299 154 300 155
rect 300 154 301 155
rect 301 154 302 155
rect 302 154 303 155
rect 303 154 304 155
rect 304 154 305 155
rect 305 154 306 155
rect 306 154 307 155
rect 336 154 337 155
rect 337 154 338 155
rect 338 154 339 155
rect 339 154 340 155
rect 340 154 341 155
rect 341 154 342 155
rect 342 154 343 155
rect 343 154 344 155
rect 344 154 345 155
rect 345 154 346 155
rect 346 154 347 155
rect 347 154 348 155
rect 375 154 376 155
rect 376 154 377 155
rect 377 154 378 155
rect 378 154 379 155
rect 379 154 380 155
rect 380 154 381 155
rect 381 154 382 155
rect 382 154 383 155
rect 383 154 384 155
rect 384 154 385 155
rect 489 154 490 155
rect 490 154 491 155
rect 491 154 492 155
rect 492 154 493 155
rect 493 154 494 155
rect 494 154 495 155
rect 495 154 496 155
rect 496 154 497 155
rect 497 154 498 155
rect 498 154 499 155
rect 499 154 500 155
rect 500 154 501 155
rect 501 154 502 155
rect 502 154 503 155
rect 503 154 504 155
rect 504 154 505 155
rect 505 154 506 155
rect 506 154 507 155
rect 507 154 508 155
rect 508 154 509 155
rect 509 154 510 155
rect 510 154 511 155
rect 511 154 512 155
rect 512 154 513 155
rect 109 153 110 154
rect 110 153 111 154
rect 111 153 112 154
rect 112 153 113 154
rect 113 153 114 154
rect 114 153 115 154
rect 115 153 116 154
rect 116 153 117 154
rect 117 153 118 154
rect 118 153 119 154
rect 208 153 209 154
rect 209 153 210 154
rect 210 153 211 154
rect 211 153 212 154
rect 212 153 213 154
rect 213 153 214 154
rect 214 153 215 154
rect 236 153 237 154
rect 237 153 238 154
rect 238 153 239 154
rect 239 153 240 154
rect 240 153 241 154
rect 241 153 242 154
rect 242 153 243 154
rect 243 153 244 154
rect 244 153 245 154
rect 245 153 246 154
rect 246 153 247 154
rect 247 153 248 154
rect 248 153 249 154
rect 278 153 279 154
rect 279 153 280 154
rect 280 153 281 154
rect 281 153 282 154
rect 282 153 283 154
rect 283 153 284 154
rect 294 153 295 154
rect 295 153 296 154
rect 296 153 297 154
rect 297 153 298 154
rect 298 153 299 154
rect 299 153 300 154
rect 300 153 301 154
rect 301 153 302 154
rect 302 153 303 154
rect 303 153 304 154
rect 304 153 305 154
rect 305 153 306 154
rect 306 153 307 154
rect 336 153 337 154
rect 337 153 338 154
rect 338 153 339 154
rect 339 153 340 154
rect 340 153 341 154
rect 341 153 342 154
rect 342 153 343 154
rect 343 153 344 154
rect 344 153 345 154
rect 345 153 346 154
rect 375 153 376 154
rect 376 153 377 154
rect 377 153 378 154
rect 378 153 379 154
rect 379 153 380 154
rect 380 153 381 154
rect 381 153 382 154
rect 382 153 383 154
rect 383 153 384 154
rect 489 153 490 154
rect 490 153 491 154
rect 491 153 492 154
rect 492 153 493 154
rect 493 153 494 154
rect 494 153 495 154
rect 495 153 496 154
rect 496 153 497 154
rect 497 153 498 154
rect 498 153 499 154
rect 499 153 500 154
rect 500 153 501 154
rect 501 153 502 154
rect 502 153 503 154
rect 503 153 504 154
rect 504 153 505 154
rect 505 153 506 154
rect 506 153 507 154
rect 507 153 508 154
rect 508 153 509 154
rect 509 153 510 154
rect 510 153 511 154
rect 109 152 110 153
rect 110 152 111 153
rect 111 152 112 153
rect 112 152 113 153
rect 113 152 114 153
rect 114 152 115 153
rect 115 152 116 153
rect 116 152 117 153
rect 117 152 118 153
rect 118 152 119 153
rect 119 152 120 153
rect 120 152 121 153
rect 208 152 209 153
rect 209 152 210 153
rect 210 152 211 153
rect 211 152 212 153
rect 212 152 213 153
rect 213 152 214 153
rect 214 152 215 153
rect 236 152 237 153
rect 237 152 238 153
rect 238 152 239 153
rect 239 152 240 153
rect 240 152 241 153
rect 241 152 242 153
rect 242 152 243 153
rect 243 152 244 153
rect 244 152 245 153
rect 245 152 246 153
rect 246 152 247 153
rect 247 152 248 153
rect 248 152 249 153
rect 276 152 277 153
rect 277 152 278 153
rect 278 152 279 153
rect 279 152 280 153
rect 280 152 281 153
rect 281 152 282 153
rect 282 152 283 153
rect 283 152 284 153
rect 294 152 295 153
rect 295 152 296 153
rect 296 152 297 153
rect 297 152 298 153
rect 298 152 299 153
rect 299 152 300 153
rect 300 152 301 153
rect 301 152 302 153
rect 302 152 303 153
rect 303 152 304 153
rect 304 152 305 153
rect 305 152 306 153
rect 306 152 307 153
rect 336 152 337 153
rect 337 152 338 153
rect 338 152 339 153
rect 339 152 340 153
rect 340 152 341 153
rect 341 152 342 153
rect 342 152 343 153
rect 343 152 344 153
rect 344 152 345 153
rect 345 152 346 153
rect 346 152 347 153
rect 347 152 348 153
rect 375 152 376 153
rect 376 152 377 153
rect 377 152 378 153
rect 378 152 379 153
rect 379 152 380 153
rect 380 152 381 153
rect 381 152 382 153
rect 382 152 383 153
rect 383 152 384 153
rect 487 152 488 153
rect 488 152 489 153
rect 489 152 490 153
rect 490 152 491 153
rect 491 152 492 153
rect 492 152 493 153
rect 493 152 494 153
rect 494 152 495 153
rect 495 152 496 153
rect 496 152 497 153
rect 497 152 498 153
rect 498 152 499 153
rect 499 152 500 153
rect 500 152 501 153
rect 501 152 502 153
rect 502 152 503 153
rect 503 152 504 153
rect 504 152 505 153
rect 505 152 506 153
rect 506 152 507 153
rect 507 152 508 153
rect 508 152 509 153
rect 509 152 510 153
rect 510 152 511 153
rect 109 151 110 152
rect 110 151 111 152
rect 111 151 112 152
rect 112 151 113 152
rect 113 151 114 152
rect 114 151 115 152
rect 115 151 116 152
rect 116 151 117 152
rect 117 151 118 152
rect 118 151 119 152
rect 119 151 120 152
rect 120 151 121 152
rect 208 151 209 152
rect 209 151 210 152
rect 210 151 211 152
rect 211 151 212 152
rect 212 151 213 152
rect 213 151 214 152
rect 214 151 215 152
rect 238 151 239 152
rect 239 151 240 152
rect 240 151 241 152
rect 241 151 242 152
rect 242 151 243 152
rect 243 151 244 152
rect 244 151 245 152
rect 245 151 246 152
rect 246 151 247 152
rect 247 151 248 152
rect 248 151 249 152
rect 276 151 277 152
rect 277 151 278 152
rect 278 151 279 152
rect 279 151 280 152
rect 280 151 281 152
rect 281 151 282 152
rect 296 151 297 152
rect 297 151 298 152
rect 298 151 299 152
rect 299 151 300 152
rect 300 151 301 152
rect 301 151 302 152
rect 302 151 303 152
rect 303 151 304 152
rect 304 151 305 152
rect 305 151 306 152
rect 306 151 307 152
rect 336 151 337 152
rect 337 151 338 152
rect 338 151 339 152
rect 339 151 340 152
rect 340 151 341 152
rect 341 151 342 152
rect 342 151 343 152
rect 343 151 344 152
rect 344 151 345 152
rect 345 151 346 152
rect 346 151 347 152
rect 347 151 348 152
rect 375 151 376 152
rect 376 151 377 152
rect 377 151 378 152
rect 378 151 379 152
rect 379 151 380 152
rect 380 151 381 152
rect 381 151 382 152
rect 487 151 488 152
rect 488 151 489 152
rect 489 151 490 152
rect 490 151 491 152
rect 491 151 492 152
rect 492 151 493 152
rect 493 151 494 152
rect 494 151 495 152
rect 495 151 496 152
rect 496 151 497 152
rect 497 151 498 152
rect 498 151 499 152
rect 499 151 500 152
rect 500 151 501 152
rect 501 151 502 152
rect 502 151 503 152
rect 503 151 504 152
rect 504 151 505 152
rect 505 151 506 152
rect 506 151 507 152
rect 507 151 508 152
rect 508 151 509 152
rect 109 150 110 151
rect 110 150 111 151
rect 111 150 112 151
rect 112 150 113 151
rect 113 150 114 151
rect 114 150 115 151
rect 115 150 116 151
rect 116 150 117 151
rect 117 150 118 151
rect 118 150 119 151
rect 119 150 120 151
rect 120 150 121 151
rect 206 150 207 151
rect 207 150 208 151
rect 208 150 209 151
rect 209 150 210 151
rect 210 150 211 151
rect 211 150 212 151
rect 212 150 213 151
rect 213 150 214 151
rect 214 150 215 151
rect 238 150 239 151
rect 239 150 240 151
rect 240 150 241 151
rect 241 150 242 151
rect 242 150 243 151
rect 243 150 244 151
rect 244 150 245 151
rect 245 150 246 151
rect 246 150 247 151
rect 247 150 248 151
rect 248 150 249 151
rect 249 150 250 151
rect 250 150 251 151
rect 276 150 277 151
rect 277 150 278 151
rect 278 150 279 151
rect 279 150 280 151
rect 280 150 281 151
rect 281 150 282 151
rect 296 150 297 151
rect 297 150 298 151
rect 298 150 299 151
rect 299 150 300 151
rect 300 150 301 151
rect 301 150 302 151
rect 302 150 303 151
rect 303 150 304 151
rect 304 150 305 151
rect 305 150 306 151
rect 306 150 307 151
rect 307 150 308 151
rect 308 150 309 151
rect 336 150 337 151
rect 337 150 338 151
rect 338 150 339 151
rect 339 150 340 151
rect 340 150 341 151
rect 341 150 342 151
rect 342 150 343 151
rect 343 150 344 151
rect 344 150 345 151
rect 345 150 346 151
rect 346 150 347 151
rect 347 150 348 151
rect 373 150 374 151
rect 374 150 375 151
rect 375 150 376 151
rect 376 150 377 151
rect 377 150 378 151
rect 378 150 379 151
rect 379 150 380 151
rect 380 150 381 151
rect 381 150 382 151
rect 409 150 410 151
rect 410 150 411 151
rect 411 150 412 151
rect 487 150 488 151
rect 488 150 489 151
rect 489 150 490 151
rect 490 150 491 151
rect 491 150 492 151
rect 492 150 493 151
rect 493 150 494 151
rect 494 150 495 151
rect 495 150 496 151
rect 496 150 497 151
rect 497 150 498 151
rect 498 150 499 151
rect 499 150 500 151
rect 500 150 501 151
rect 501 150 502 151
rect 502 150 503 151
rect 503 150 504 151
rect 504 150 505 151
rect 505 150 506 151
rect 506 150 507 151
rect 507 150 508 151
rect 508 150 509 151
rect 111 149 112 150
rect 112 149 113 150
rect 113 149 114 150
rect 114 149 115 150
rect 115 149 116 150
rect 116 149 117 150
rect 117 149 118 150
rect 118 149 119 150
rect 119 149 120 150
rect 120 149 121 150
rect 206 149 207 150
rect 207 149 208 150
rect 208 149 209 150
rect 209 149 210 150
rect 210 149 211 150
rect 211 149 212 150
rect 212 149 213 150
rect 238 149 239 150
rect 239 149 240 150
rect 240 149 241 150
rect 241 149 242 150
rect 242 149 243 150
rect 243 149 244 150
rect 244 149 245 150
rect 245 149 246 150
rect 246 149 247 150
rect 247 149 248 150
rect 248 149 249 150
rect 249 149 250 150
rect 250 149 251 150
rect 276 149 277 150
rect 277 149 278 150
rect 278 149 279 150
rect 279 149 280 150
rect 280 149 281 150
rect 281 149 282 150
rect 296 149 297 150
rect 297 149 298 150
rect 298 149 299 150
rect 299 149 300 150
rect 300 149 301 150
rect 301 149 302 150
rect 302 149 303 150
rect 303 149 304 150
rect 304 149 305 150
rect 305 149 306 150
rect 306 149 307 150
rect 307 149 308 150
rect 308 149 309 150
rect 336 149 337 150
rect 337 149 338 150
rect 338 149 339 150
rect 339 149 340 150
rect 340 149 341 150
rect 341 149 342 150
rect 342 149 343 150
rect 343 149 344 150
rect 344 149 345 150
rect 345 149 346 150
rect 373 149 374 150
rect 374 149 375 150
rect 375 149 376 150
rect 376 149 377 150
rect 377 149 378 150
rect 378 149 379 150
rect 379 149 380 150
rect 380 149 381 150
rect 381 149 382 150
rect 409 149 410 150
rect 410 149 411 150
rect 411 149 412 150
rect 487 149 488 150
rect 488 149 489 150
rect 489 149 490 150
rect 490 149 491 150
rect 491 149 492 150
rect 492 149 493 150
rect 493 149 494 150
rect 494 149 495 150
rect 495 149 496 150
rect 496 149 497 150
rect 497 149 498 150
rect 498 149 499 150
rect 499 149 500 150
rect 500 149 501 150
rect 501 149 502 150
rect 502 149 503 150
rect 503 149 504 150
rect 504 149 505 150
rect 505 149 506 150
rect 506 149 507 150
rect 111 148 112 149
rect 112 148 113 149
rect 113 148 114 149
rect 114 148 115 149
rect 115 148 116 149
rect 116 148 117 149
rect 117 148 118 149
rect 118 148 119 149
rect 119 148 120 149
rect 120 148 121 149
rect 121 148 122 149
rect 122 148 123 149
rect 206 148 207 149
rect 207 148 208 149
rect 208 148 209 149
rect 209 148 210 149
rect 210 148 211 149
rect 211 148 212 149
rect 212 148 213 149
rect 238 148 239 149
rect 239 148 240 149
rect 240 148 241 149
rect 241 148 242 149
rect 242 148 243 149
rect 243 148 244 149
rect 244 148 245 149
rect 245 148 246 149
rect 246 148 247 149
rect 247 148 248 149
rect 248 148 249 149
rect 249 148 250 149
rect 250 148 251 149
rect 251 148 252 149
rect 276 148 277 149
rect 277 148 278 149
rect 278 148 279 149
rect 279 148 280 149
rect 280 148 281 149
rect 281 148 282 149
rect 296 148 297 149
rect 297 148 298 149
rect 298 148 299 149
rect 299 148 300 149
rect 300 148 301 149
rect 301 148 302 149
rect 302 148 303 149
rect 303 148 304 149
rect 304 148 305 149
rect 305 148 306 149
rect 306 148 307 149
rect 307 148 308 149
rect 308 148 309 149
rect 336 148 337 149
rect 337 148 338 149
rect 338 148 339 149
rect 339 148 340 149
rect 340 148 341 149
rect 341 148 342 149
rect 342 148 343 149
rect 343 148 344 149
rect 344 148 345 149
rect 345 148 346 149
rect 371 148 372 149
rect 372 148 373 149
rect 373 148 374 149
rect 374 148 375 149
rect 375 148 376 149
rect 376 148 377 149
rect 377 148 378 149
rect 378 148 379 149
rect 379 148 380 149
rect 380 148 381 149
rect 381 148 382 149
rect 407 148 408 149
rect 408 148 409 149
rect 409 148 410 149
rect 410 148 411 149
rect 411 148 412 149
rect 486 148 487 149
rect 487 148 488 149
rect 488 148 489 149
rect 489 148 490 149
rect 490 148 491 149
rect 491 148 492 149
rect 492 148 493 149
rect 493 148 494 149
rect 494 148 495 149
rect 495 148 496 149
rect 496 148 497 149
rect 497 148 498 149
rect 498 148 499 149
rect 499 148 500 149
rect 500 148 501 149
rect 501 148 502 149
rect 502 148 503 149
rect 503 148 504 149
rect 504 148 505 149
rect 505 148 506 149
rect 506 148 507 149
rect 111 147 112 148
rect 112 147 113 148
rect 113 147 114 148
rect 114 147 115 148
rect 115 147 116 148
rect 116 147 117 148
rect 117 147 118 148
rect 118 147 119 148
rect 119 147 120 148
rect 120 147 121 148
rect 121 147 122 148
rect 122 147 123 148
rect 206 147 207 148
rect 207 147 208 148
rect 208 147 209 148
rect 209 147 210 148
rect 210 147 211 148
rect 211 147 212 148
rect 212 147 213 148
rect 238 147 239 148
rect 239 147 240 148
rect 240 147 241 148
rect 241 147 242 148
rect 242 147 243 148
rect 243 147 244 148
rect 244 147 245 148
rect 245 147 246 148
rect 246 147 247 148
rect 247 147 248 148
rect 248 147 249 148
rect 249 147 250 148
rect 250 147 251 148
rect 251 147 252 148
rect 276 147 277 148
rect 277 147 278 148
rect 278 147 279 148
rect 279 147 280 148
rect 296 147 297 148
rect 297 147 298 148
rect 298 147 299 148
rect 299 147 300 148
rect 300 147 301 148
rect 301 147 302 148
rect 302 147 303 148
rect 303 147 304 148
rect 304 147 305 148
rect 305 147 306 148
rect 306 147 307 148
rect 307 147 308 148
rect 308 147 309 148
rect 336 147 337 148
rect 337 147 338 148
rect 338 147 339 148
rect 339 147 340 148
rect 340 147 341 148
rect 341 147 342 148
rect 342 147 343 148
rect 343 147 344 148
rect 344 147 345 148
rect 345 147 346 148
rect 371 147 372 148
rect 372 147 373 148
rect 373 147 374 148
rect 374 147 375 148
rect 375 147 376 148
rect 376 147 377 148
rect 377 147 378 148
rect 407 147 408 148
rect 408 147 409 148
rect 409 147 410 148
rect 410 147 411 148
rect 411 147 412 148
rect 486 147 487 148
rect 487 147 488 148
rect 488 147 489 148
rect 489 147 490 148
rect 490 147 491 148
rect 491 147 492 148
rect 492 147 493 148
rect 493 147 494 148
rect 494 147 495 148
rect 495 147 496 148
rect 496 147 497 148
rect 497 147 498 148
rect 498 147 499 148
rect 499 147 500 148
rect 500 147 501 148
rect 501 147 502 148
rect 502 147 503 148
rect 503 147 504 148
rect 504 147 505 148
rect 111 146 112 147
rect 112 146 113 147
rect 113 146 114 147
rect 114 146 115 147
rect 115 146 116 147
rect 116 146 117 147
rect 117 146 118 147
rect 118 146 119 147
rect 119 146 120 147
rect 120 146 121 147
rect 121 146 122 147
rect 122 146 123 147
rect 206 146 207 147
rect 207 146 208 147
rect 208 146 209 147
rect 209 146 210 147
rect 210 146 211 147
rect 211 146 212 147
rect 212 146 213 147
rect 238 146 239 147
rect 239 146 240 147
rect 240 146 241 147
rect 241 146 242 147
rect 242 146 243 147
rect 243 146 244 147
rect 244 146 245 147
rect 245 146 246 147
rect 246 146 247 147
rect 247 146 248 147
rect 248 146 249 147
rect 249 146 250 147
rect 250 146 251 147
rect 251 146 252 147
rect 274 146 275 147
rect 275 146 276 147
rect 276 146 277 147
rect 277 146 278 147
rect 278 146 279 147
rect 279 146 280 147
rect 296 146 297 147
rect 297 146 298 147
rect 298 146 299 147
rect 299 146 300 147
rect 300 146 301 147
rect 301 146 302 147
rect 302 146 303 147
rect 303 146 304 147
rect 304 146 305 147
rect 305 146 306 147
rect 306 146 307 147
rect 307 146 308 147
rect 308 146 309 147
rect 309 146 310 147
rect 336 146 337 147
rect 337 146 338 147
rect 338 146 339 147
rect 339 146 340 147
rect 340 146 341 147
rect 341 146 342 147
rect 342 146 343 147
rect 343 146 344 147
rect 344 146 345 147
rect 345 146 346 147
rect 369 146 370 147
rect 370 146 371 147
rect 371 146 372 147
rect 372 146 373 147
rect 373 146 374 147
rect 374 146 375 147
rect 375 146 376 147
rect 376 146 377 147
rect 377 146 378 147
rect 407 146 408 147
rect 408 146 409 147
rect 409 146 410 147
rect 410 146 411 147
rect 411 146 412 147
rect 484 146 485 147
rect 485 146 486 147
rect 486 146 487 147
rect 487 146 488 147
rect 488 146 489 147
rect 489 146 490 147
rect 490 146 491 147
rect 491 146 492 147
rect 492 146 493 147
rect 493 146 494 147
rect 494 146 495 147
rect 495 146 496 147
rect 496 146 497 147
rect 497 146 498 147
rect 498 146 499 147
rect 499 146 500 147
rect 500 146 501 147
rect 501 146 502 147
rect 502 146 503 147
rect 503 146 504 147
rect 504 146 505 147
rect 113 145 114 146
rect 114 145 115 146
rect 115 145 116 146
rect 116 145 117 146
rect 117 145 118 146
rect 118 145 119 146
rect 119 145 120 146
rect 120 145 121 146
rect 121 145 122 146
rect 122 145 123 146
rect 206 145 207 146
rect 207 145 208 146
rect 208 145 209 146
rect 209 145 210 146
rect 210 145 211 146
rect 240 145 241 146
rect 241 145 242 146
rect 242 145 243 146
rect 243 145 244 146
rect 244 145 245 146
rect 245 145 246 146
rect 246 145 247 146
rect 247 145 248 146
rect 248 145 249 146
rect 249 145 250 146
rect 250 145 251 146
rect 251 145 252 146
rect 274 145 275 146
rect 275 145 276 146
rect 276 145 277 146
rect 277 145 278 146
rect 278 145 279 146
rect 279 145 280 146
rect 298 145 299 146
rect 299 145 300 146
rect 300 145 301 146
rect 301 145 302 146
rect 302 145 303 146
rect 303 145 304 146
rect 304 145 305 146
rect 305 145 306 146
rect 306 145 307 146
rect 307 145 308 146
rect 308 145 309 146
rect 309 145 310 146
rect 336 145 337 146
rect 337 145 338 146
rect 338 145 339 146
rect 339 145 340 146
rect 340 145 341 146
rect 341 145 342 146
rect 342 145 343 146
rect 343 145 344 146
rect 344 145 345 146
rect 345 145 346 146
rect 369 145 370 146
rect 370 145 371 146
rect 371 145 372 146
rect 372 145 373 146
rect 373 145 374 146
rect 374 145 375 146
rect 375 145 376 146
rect 376 145 377 146
rect 377 145 378 146
rect 407 145 408 146
rect 408 145 409 146
rect 409 145 410 146
rect 410 145 411 146
rect 411 145 412 146
rect 484 145 485 146
rect 485 145 486 146
rect 486 145 487 146
rect 487 145 488 146
rect 488 145 489 146
rect 489 145 490 146
rect 490 145 491 146
rect 491 145 492 146
rect 492 145 493 146
rect 493 145 494 146
rect 494 145 495 146
rect 495 145 496 146
rect 496 145 497 146
rect 497 145 498 146
rect 498 145 499 146
rect 499 145 500 146
rect 500 145 501 146
rect 501 145 502 146
rect 502 145 503 146
rect 113 144 114 145
rect 114 144 115 145
rect 115 144 116 145
rect 116 144 117 145
rect 117 144 118 145
rect 118 144 119 145
rect 119 144 120 145
rect 120 144 121 145
rect 121 144 122 145
rect 122 144 123 145
rect 123 144 124 145
rect 124 144 125 145
rect 203 144 204 145
rect 204 144 205 145
rect 205 144 206 145
rect 206 144 207 145
rect 207 144 208 145
rect 208 144 209 145
rect 209 144 210 145
rect 210 144 211 145
rect 211 144 212 145
rect 212 144 213 145
rect 238 144 239 145
rect 239 144 240 145
rect 240 144 241 145
rect 241 144 242 145
rect 242 144 243 145
rect 243 144 244 145
rect 244 144 245 145
rect 245 144 246 145
rect 246 144 247 145
rect 247 144 248 145
rect 248 144 249 145
rect 249 144 250 145
rect 250 144 251 145
rect 251 144 252 145
rect 252 144 253 145
rect 253 144 254 145
rect 274 144 275 145
rect 275 144 276 145
rect 276 144 277 145
rect 277 144 278 145
rect 278 144 279 145
rect 279 144 280 145
rect 298 144 299 145
rect 299 144 300 145
rect 300 144 301 145
rect 301 144 302 145
rect 302 144 303 145
rect 303 144 304 145
rect 304 144 305 145
rect 305 144 306 145
rect 306 144 307 145
rect 307 144 308 145
rect 308 144 309 145
rect 309 144 310 145
rect 336 144 337 145
rect 337 144 338 145
rect 338 144 339 145
rect 339 144 340 145
rect 340 144 341 145
rect 341 144 342 145
rect 342 144 343 145
rect 343 144 344 145
rect 344 144 345 145
rect 345 144 346 145
rect 346 144 347 145
rect 347 144 348 145
rect 369 144 370 145
rect 370 144 371 145
rect 371 144 372 145
rect 372 144 373 145
rect 373 144 374 145
rect 374 144 375 145
rect 375 144 376 145
rect 376 144 377 145
rect 377 144 378 145
rect 405 144 406 145
rect 406 144 407 145
rect 407 144 408 145
rect 408 144 409 145
rect 409 144 410 145
rect 410 144 411 145
rect 411 144 412 145
rect 482 144 483 145
rect 483 144 484 145
rect 484 144 485 145
rect 485 144 486 145
rect 486 144 487 145
rect 487 144 488 145
rect 488 144 489 145
rect 489 144 490 145
rect 490 144 491 145
rect 491 144 492 145
rect 492 144 493 145
rect 493 144 494 145
rect 494 144 495 145
rect 495 144 496 145
rect 496 144 497 145
rect 497 144 498 145
rect 498 144 499 145
rect 499 144 500 145
rect 500 144 501 145
rect 501 144 502 145
rect 502 144 503 145
rect 113 143 114 144
rect 114 143 115 144
rect 115 143 116 144
rect 116 143 117 144
rect 117 143 118 144
rect 118 143 119 144
rect 119 143 120 144
rect 120 143 121 144
rect 121 143 122 144
rect 122 143 123 144
rect 123 143 124 144
rect 124 143 125 144
rect 203 143 204 144
rect 204 143 205 144
rect 205 143 206 144
rect 206 143 207 144
rect 207 143 208 144
rect 208 143 209 144
rect 209 143 210 144
rect 210 143 211 144
rect 211 143 212 144
rect 212 143 213 144
rect 238 143 239 144
rect 239 143 240 144
rect 240 143 241 144
rect 241 143 242 144
rect 242 143 243 144
rect 243 143 244 144
rect 244 143 245 144
rect 245 143 246 144
rect 246 143 247 144
rect 247 143 248 144
rect 248 143 249 144
rect 249 143 250 144
rect 250 143 251 144
rect 251 143 252 144
rect 252 143 253 144
rect 253 143 254 144
rect 274 143 275 144
rect 275 143 276 144
rect 276 143 277 144
rect 277 143 278 144
rect 278 143 279 144
rect 279 143 280 144
rect 298 143 299 144
rect 299 143 300 144
rect 300 143 301 144
rect 301 143 302 144
rect 302 143 303 144
rect 303 143 304 144
rect 304 143 305 144
rect 305 143 306 144
rect 306 143 307 144
rect 307 143 308 144
rect 308 143 309 144
rect 309 143 310 144
rect 336 143 337 144
rect 337 143 338 144
rect 338 143 339 144
rect 339 143 340 144
rect 340 143 341 144
rect 341 143 342 144
rect 342 143 343 144
rect 343 143 344 144
rect 344 143 345 144
rect 345 143 346 144
rect 346 143 347 144
rect 347 143 348 144
rect 369 143 370 144
rect 370 143 371 144
rect 371 143 372 144
rect 372 143 373 144
rect 373 143 374 144
rect 405 143 406 144
rect 406 143 407 144
rect 407 143 408 144
rect 408 143 409 144
rect 409 143 410 144
rect 410 143 411 144
rect 411 143 412 144
rect 482 143 483 144
rect 483 143 484 144
rect 484 143 485 144
rect 485 143 486 144
rect 486 143 487 144
rect 487 143 488 144
rect 488 143 489 144
rect 489 143 490 144
rect 490 143 491 144
rect 491 143 492 144
rect 492 143 493 144
rect 493 143 494 144
rect 494 143 495 144
rect 495 143 496 144
rect 496 143 497 144
rect 497 143 498 144
rect 498 143 499 144
rect 499 143 500 144
rect 500 143 501 144
rect 501 143 502 144
rect 113 142 114 143
rect 114 142 115 143
rect 115 142 116 143
rect 116 142 117 143
rect 117 142 118 143
rect 118 142 119 143
rect 119 142 120 143
rect 120 142 121 143
rect 121 142 122 143
rect 122 142 123 143
rect 123 142 124 143
rect 124 142 125 143
rect 125 142 126 143
rect 126 142 127 143
rect 199 142 200 143
rect 200 142 201 143
rect 201 142 202 143
rect 202 142 203 143
rect 203 142 204 143
rect 204 142 205 143
rect 205 142 206 143
rect 206 142 207 143
rect 207 142 208 143
rect 208 142 209 143
rect 209 142 210 143
rect 210 142 211 143
rect 211 142 212 143
rect 212 142 213 143
rect 213 142 214 143
rect 214 142 215 143
rect 236 142 237 143
rect 237 142 238 143
rect 238 142 239 143
rect 239 142 240 143
rect 240 142 241 143
rect 241 142 242 143
rect 242 142 243 143
rect 243 142 244 143
rect 244 142 245 143
rect 245 142 246 143
rect 246 142 247 143
rect 247 142 248 143
rect 248 142 249 143
rect 249 142 250 143
rect 250 142 251 143
rect 251 142 252 143
rect 252 142 253 143
rect 253 142 254 143
rect 254 142 255 143
rect 255 142 256 143
rect 274 142 275 143
rect 275 142 276 143
rect 276 142 277 143
rect 277 142 278 143
rect 278 142 279 143
rect 279 142 280 143
rect 298 142 299 143
rect 299 142 300 143
rect 300 142 301 143
rect 301 142 302 143
rect 302 142 303 143
rect 303 142 304 143
rect 304 142 305 143
rect 305 142 306 143
rect 306 142 307 143
rect 307 142 308 143
rect 308 142 309 143
rect 309 142 310 143
rect 336 142 337 143
rect 337 142 338 143
rect 338 142 339 143
rect 339 142 340 143
rect 340 142 341 143
rect 341 142 342 143
rect 342 142 343 143
rect 343 142 344 143
rect 344 142 345 143
rect 345 142 346 143
rect 346 142 347 143
rect 347 142 348 143
rect 366 142 367 143
rect 367 142 368 143
rect 368 142 369 143
rect 369 142 370 143
rect 370 142 371 143
rect 371 142 372 143
rect 372 142 373 143
rect 373 142 374 143
rect 403 142 404 143
rect 404 142 405 143
rect 405 142 406 143
rect 406 142 407 143
rect 407 142 408 143
rect 408 142 409 143
rect 409 142 410 143
rect 410 142 411 143
rect 411 142 412 143
rect 480 142 481 143
rect 481 142 482 143
rect 482 142 483 143
rect 483 142 484 143
rect 484 142 485 143
rect 485 142 486 143
rect 486 142 487 143
rect 487 142 488 143
rect 488 142 489 143
rect 489 142 490 143
rect 490 142 491 143
rect 491 142 492 143
rect 492 142 493 143
rect 493 142 494 143
rect 494 142 495 143
rect 495 142 496 143
rect 496 142 497 143
rect 497 142 498 143
rect 498 142 499 143
rect 499 142 500 143
rect 500 142 501 143
rect 501 142 502 143
rect 115 141 116 142
rect 116 141 117 142
rect 117 141 118 142
rect 118 141 119 142
rect 119 141 120 142
rect 120 141 121 142
rect 121 141 122 142
rect 122 141 123 142
rect 123 141 124 142
rect 124 141 125 142
rect 125 141 126 142
rect 126 141 127 142
rect 199 141 200 142
rect 200 141 201 142
rect 201 141 202 142
rect 202 141 203 142
rect 203 141 204 142
rect 204 141 205 142
rect 205 141 206 142
rect 206 141 207 142
rect 207 141 208 142
rect 208 141 209 142
rect 209 141 210 142
rect 210 141 211 142
rect 211 141 212 142
rect 212 141 213 142
rect 213 141 214 142
rect 214 141 215 142
rect 236 141 237 142
rect 237 141 238 142
rect 238 141 239 142
rect 239 141 240 142
rect 240 141 241 142
rect 241 141 242 142
rect 242 141 243 142
rect 243 141 244 142
rect 244 141 245 142
rect 245 141 246 142
rect 246 141 247 142
rect 247 141 248 142
rect 248 141 249 142
rect 249 141 250 142
rect 250 141 251 142
rect 251 141 252 142
rect 252 141 253 142
rect 253 141 254 142
rect 254 141 255 142
rect 255 141 256 142
rect 274 141 275 142
rect 275 141 276 142
rect 276 141 277 142
rect 277 141 278 142
rect 278 141 279 142
rect 300 141 301 142
rect 301 141 302 142
rect 302 141 303 142
rect 303 141 304 142
rect 304 141 305 142
rect 305 141 306 142
rect 306 141 307 142
rect 307 141 308 142
rect 308 141 309 142
rect 309 141 310 142
rect 336 141 337 142
rect 337 141 338 142
rect 338 141 339 142
rect 339 141 340 142
rect 340 141 341 142
rect 341 141 342 142
rect 342 141 343 142
rect 343 141 344 142
rect 344 141 345 142
rect 345 141 346 142
rect 366 141 367 142
rect 367 141 368 142
rect 368 141 369 142
rect 369 141 370 142
rect 370 141 371 142
rect 371 141 372 142
rect 372 141 373 142
rect 373 141 374 142
rect 403 141 404 142
rect 404 141 405 142
rect 405 141 406 142
rect 406 141 407 142
rect 407 141 408 142
rect 408 141 409 142
rect 409 141 410 142
rect 410 141 411 142
rect 411 141 412 142
rect 480 141 481 142
rect 481 141 482 142
rect 482 141 483 142
rect 483 141 484 142
rect 484 141 485 142
rect 485 141 486 142
rect 486 141 487 142
rect 487 141 488 142
rect 488 141 489 142
rect 489 141 490 142
rect 490 141 491 142
rect 491 141 492 142
rect 492 141 493 142
rect 493 141 494 142
rect 494 141 495 142
rect 495 141 496 142
rect 496 141 497 142
rect 497 141 498 142
rect 498 141 499 142
rect 499 141 500 142
rect 500 141 501 142
rect 501 141 502 142
rect 115 140 116 141
rect 116 140 117 141
rect 117 140 118 141
rect 118 140 119 141
rect 119 140 120 141
rect 120 140 121 141
rect 121 140 122 141
rect 122 140 123 141
rect 123 140 124 141
rect 124 140 125 141
rect 125 140 126 141
rect 126 140 127 141
rect 197 140 198 141
rect 198 140 199 141
rect 199 140 200 141
rect 200 140 201 141
rect 201 140 202 141
rect 202 140 203 141
rect 203 140 204 141
rect 204 140 205 141
rect 205 140 206 141
rect 206 140 207 141
rect 207 140 208 141
rect 208 140 209 141
rect 209 140 210 141
rect 210 140 211 141
rect 211 140 212 141
rect 212 140 213 141
rect 213 140 214 141
rect 214 140 215 141
rect 215 140 216 141
rect 216 140 217 141
rect 217 140 218 141
rect 218 140 219 141
rect 233 140 234 141
rect 234 140 235 141
rect 235 140 236 141
rect 236 140 237 141
rect 237 140 238 141
rect 238 140 239 141
rect 239 140 240 141
rect 240 140 241 141
rect 241 140 242 141
rect 242 140 243 141
rect 243 140 244 141
rect 244 140 245 141
rect 245 140 246 141
rect 246 140 247 141
rect 247 140 248 141
rect 248 140 249 141
rect 249 140 250 141
rect 250 140 251 141
rect 251 140 252 141
rect 252 140 253 141
rect 253 140 254 141
rect 254 140 255 141
rect 255 140 256 141
rect 256 140 257 141
rect 257 140 258 141
rect 258 140 259 141
rect 259 140 260 141
rect 272 140 273 141
rect 273 140 274 141
rect 274 140 275 141
rect 275 140 276 141
rect 276 140 277 141
rect 277 140 278 141
rect 278 140 279 141
rect 300 140 301 141
rect 301 140 302 141
rect 302 140 303 141
rect 303 140 304 141
rect 304 140 305 141
rect 305 140 306 141
rect 306 140 307 141
rect 307 140 308 141
rect 308 140 309 141
rect 309 140 310 141
rect 310 140 311 141
rect 311 140 312 141
rect 336 140 337 141
rect 337 140 338 141
rect 338 140 339 141
rect 339 140 340 141
rect 340 140 341 141
rect 341 140 342 141
rect 342 140 343 141
rect 343 140 344 141
rect 344 140 345 141
rect 345 140 346 141
rect 366 140 367 141
rect 367 140 368 141
rect 368 140 369 141
rect 369 140 370 141
rect 370 140 371 141
rect 371 140 372 141
rect 372 140 373 141
rect 373 140 374 141
rect 374 140 375 141
rect 375 140 376 141
rect 376 140 377 141
rect 377 140 378 141
rect 379 140 380 141
rect 380 140 381 141
rect 381 140 382 141
rect 382 140 383 141
rect 383 140 384 141
rect 384 140 385 141
rect 385 140 386 141
rect 386 140 387 141
rect 387 140 388 141
rect 388 140 389 141
rect 390 140 391 141
rect 391 140 392 141
rect 392 140 393 141
rect 393 140 394 141
rect 394 140 395 141
rect 395 140 396 141
rect 396 140 397 141
rect 397 140 398 141
rect 398 140 399 141
rect 399 140 400 141
rect 400 140 401 141
rect 401 140 402 141
rect 402 140 403 141
rect 403 140 404 141
rect 404 140 405 141
rect 405 140 406 141
rect 406 140 407 141
rect 407 140 408 141
rect 408 140 409 141
rect 409 140 410 141
rect 410 140 411 141
rect 411 140 412 141
rect 478 140 479 141
rect 479 140 480 141
rect 480 140 481 141
rect 481 140 482 141
rect 482 140 483 141
rect 483 140 484 141
rect 484 140 485 141
rect 485 140 486 141
rect 486 140 487 141
rect 487 140 488 141
rect 488 140 489 141
rect 489 140 490 141
rect 490 140 491 141
rect 491 140 492 141
rect 492 140 493 141
rect 493 140 494 141
rect 494 140 495 141
rect 495 140 496 141
rect 496 140 497 141
rect 497 140 498 141
rect 498 140 499 141
rect 499 140 500 141
rect 500 140 501 141
rect 501 140 502 141
rect 115 139 116 140
rect 116 139 117 140
rect 117 139 118 140
rect 118 139 119 140
rect 119 139 120 140
rect 120 139 121 140
rect 121 139 122 140
rect 122 139 123 140
rect 123 139 124 140
rect 124 139 125 140
rect 125 139 126 140
rect 126 139 127 140
rect 197 139 198 140
rect 198 139 199 140
rect 199 139 200 140
rect 200 139 201 140
rect 201 139 202 140
rect 202 139 203 140
rect 203 139 204 140
rect 204 139 205 140
rect 205 139 206 140
rect 206 139 207 140
rect 207 139 208 140
rect 208 139 209 140
rect 209 139 210 140
rect 210 139 211 140
rect 211 139 212 140
rect 212 139 213 140
rect 213 139 214 140
rect 214 139 215 140
rect 215 139 216 140
rect 216 139 217 140
rect 217 139 218 140
rect 218 139 219 140
rect 233 139 234 140
rect 234 139 235 140
rect 235 139 236 140
rect 236 139 237 140
rect 237 139 238 140
rect 238 139 239 140
rect 239 139 240 140
rect 240 139 241 140
rect 241 139 242 140
rect 242 139 243 140
rect 243 139 244 140
rect 244 139 245 140
rect 245 139 246 140
rect 246 139 247 140
rect 247 139 248 140
rect 248 139 249 140
rect 249 139 250 140
rect 250 139 251 140
rect 251 139 252 140
rect 252 139 253 140
rect 253 139 254 140
rect 254 139 255 140
rect 255 139 256 140
rect 256 139 257 140
rect 257 139 258 140
rect 258 139 259 140
rect 259 139 260 140
rect 272 139 273 140
rect 273 139 274 140
rect 274 139 275 140
rect 275 139 276 140
rect 276 139 277 140
rect 277 139 278 140
rect 278 139 279 140
rect 300 139 301 140
rect 301 139 302 140
rect 302 139 303 140
rect 303 139 304 140
rect 304 139 305 140
rect 305 139 306 140
rect 306 139 307 140
rect 307 139 308 140
rect 308 139 309 140
rect 309 139 310 140
rect 310 139 311 140
rect 311 139 312 140
rect 336 139 337 140
rect 337 139 338 140
rect 338 139 339 140
rect 339 139 340 140
rect 340 139 341 140
rect 341 139 342 140
rect 342 139 343 140
rect 343 139 344 140
rect 344 139 345 140
rect 345 139 346 140
rect 366 139 367 140
rect 367 139 368 140
rect 368 139 369 140
rect 369 139 370 140
rect 370 139 371 140
rect 371 139 372 140
rect 372 139 373 140
rect 373 139 374 140
rect 374 139 375 140
rect 375 139 376 140
rect 376 139 377 140
rect 377 139 378 140
rect 379 139 380 140
rect 380 139 381 140
rect 381 139 382 140
rect 382 139 383 140
rect 383 139 384 140
rect 384 139 385 140
rect 385 139 386 140
rect 386 139 387 140
rect 387 139 388 140
rect 388 139 389 140
rect 390 139 391 140
rect 391 139 392 140
rect 392 139 393 140
rect 393 139 394 140
rect 394 139 395 140
rect 395 139 396 140
rect 396 139 397 140
rect 397 139 398 140
rect 398 139 399 140
rect 399 139 400 140
rect 400 139 401 140
rect 401 139 402 140
rect 402 139 403 140
rect 403 139 404 140
rect 404 139 405 140
rect 405 139 406 140
rect 406 139 407 140
rect 407 139 408 140
rect 408 139 409 140
rect 409 139 410 140
rect 478 139 479 140
rect 479 139 480 140
rect 480 139 481 140
rect 481 139 482 140
rect 482 139 483 140
rect 483 139 484 140
rect 484 139 485 140
rect 485 139 486 140
rect 486 139 487 140
rect 487 139 488 140
rect 488 139 489 140
rect 489 139 490 140
rect 490 139 491 140
rect 491 139 492 140
rect 492 139 493 140
rect 493 139 494 140
rect 494 139 495 140
rect 495 139 496 140
rect 496 139 497 140
rect 497 139 498 140
rect 115 138 116 139
rect 116 138 117 139
rect 117 138 118 139
rect 118 138 119 139
rect 119 138 120 139
rect 120 138 121 139
rect 121 138 122 139
rect 122 138 123 139
rect 123 138 124 139
rect 124 138 125 139
rect 125 138 126 139
rect 126 138 127 139
rect 127 138 128 139
rect 128 138 129 139
rect 197 138 198 139
rect 198 138 199 139
rect 199 138 200 139
rect 200 138 201 139
rect 201 138 202 139
rect 202 138 203 139
rect 203 138 204 139
rect 204 138 205 139
rect 205 138 206 139
rect 206 138 207 139
rect 207 138 208 139
rect 208 138 209 139
rect 209 138 210 139
rect 210 138 211 139
rect 211 138 212 139
rect 212 138 213 139
rect 213 138 214 139
rect 214 138 215 139
rect 215 138 216 139
rect 216 138 217 139
rect 217 138 218 139
rect 218 138 219 139
rect 233 138 234 139
rect 234 138 235 139
rect 235 138 236 139
rect 236 138 237 139
rect 237 138 238 139
rect 238 138 239 139
rect 239 138 240 139
rect 240 138 241 139
rect 241 138 242 139
rect 242 138 243 139
rect 243 138 244 139
rect 244 138 245 139
rect 245 138 246 139
rect 246 138 247 139
rect 247 138 248 139
rect 248 138 249 139
rect 249 138 250 139
rect 250 138 251 139
rect 251 138 252 139
rect 252 138 253 139
rect 253 138 254 139
rect 254 138 255 139
rect 255 138 256 139
rect 256 138 257 139
rect 257 138 258 139
rect 258 138 259 139
rect 259 138 260 139
rect 272 138 273 139
rect 273 138 274 139
rect 274 138 275 139
rect 275 138 276 139
rect 276 138 277 139
rect 277 138 278 139
rect 278 138 279 139
rect 300 138 301 139
rect 301 138 302 139
rect 302 138 303 139
rect 303 138 304 139
rect 304 138 305 139
rect 305 138 306 139
rect 306 138 307 139
rect 307 138 308 139
rect 308 138 309 139
rect 309 138 310 139
rect 310 138 311 139
rect 311 138 312 139
rect 336 138 337 139
rect 337 138 338 139
rect 338 138 339 139
rect 339 138 340 139
rect 340 138 341 139
rect 341 138 342 139
rect 342 138 343 139
rect 343 138 344 139
rect 344 138 345 139
rect 345 138 346 139
rect 346 138 347 139
rect 347 138 348 139
rect 364 138 365 139
rect 365 138 366 139
rect 366 138 367 139
rect 367 138 368 139
rect 368 138 369 139
rect 369 138 370 139
rect 370 138 371 139
rect 371 138 372 139
rect 372 138 373 139
rect 373 138 374 139
rect 374 138 375 139
rect 375 138 376 139
rect 376 138 377 139
rect 377 138 378 139
rect 378 138 379 139
rect 379 138 380 139
rect 380 138 381 139
rect 381 138 382 139
rect 382 138 383 139
rect 383 138 384 139
rect 384 138 385 139
rect 385 138 386 139
rect 386 138 387 139
rect 387 138 388 139
rect 388 138 389 139
rect 389 138 390 139
rect 390 138 391 139
rect 391 138 392 139
rect 392 138 393 139
rect 393 138 394 139
rect 394 138 395 139
rect 395 138 396 139
rect 396 138 397 139
rect 397 138 398 139
rect 398 138 399 139
rect 399 138 400 139
rect 400 138 401 139
rect 401 138 402 139
rect 402 138 403 139
rect 403 138 404 139
rect 404 138 405 139
rect 405 138 406 139
rect 406 138 407 139
rect 407 138 408 139
rect 408 138 409 139
rect 409 138 410 139
rect 476 138 477 139
rect 477 138 478 139
rect 478 138 479 139
rect 479 138 480 139
rect 480 138 481 139
rect 481 138 482 139
rect 482 138 483 139
rect 483 138 484 139
rect 484 138 485 139
rect 485 138 486 139
rect 486 138 487 139
rect 487 138 488 139
rect 488 138 489 139
rect 489 138 490 139
rect 490 138 491 139
rect 491 138 492 139
rect 492 138 493 139
rect 493 138 494 139
rect 494 138 495 139
rect 495 138 496 139
rect 496 138 497 139
rect 497 138 498 139
rect 117 137 118 138
rect 118 137 119 138
rect 119 137 120 138
rect 120 137 121 138
rect 121 137 122 138
rect 122 137 123 138
rect 123 137 124 138
rect 124 137 125 138
rect 125 137 126 138
rect 126 137 127 138
rect 127 137 128 138
rect 128 137 129 138
rect 272 137 273 138
rect 273 137 274 138
rect 274 137 275 138
rect 275 137 276 138
rect 276 137 277 138
rect 277 137 278 138
rect 278 137 279 138
rect 300 137 301 138
rect 301 137 302 138
rect 302 137 303 138
rect 303 137 304 138
rect 304 137 305 138
rect 305 137 306 138
rect 306 137 307 138
rect 307 137 308 138
rect 308 137 309 138
rect 309 137 310 138
rect 310 137 311 138
rect 311 137 312 138
rect 336 137 337 138
rect 337 137 338 138
rect 338 137 339 138
rect 339 137 340 138
rect 340 137 341 138
rect 341 137 342 138
rect 342 137 343 138
rect 343 137 344 138
rect 344 137 345 138
rect 345 137 346 138
rect 346 137 347 138
rect 347 137 348 138
rect 364 137 365 138
rect 365 137 366 138
rect 366 137 367 138
rect 367 137 368 138
rect 368 137 369 138
rect 369 137 370 138
rect 370 137 371 138
rect 371 137 372 138
rect 372 137 373 138
rect 373 137 374 138
rect 374 137 375 138
rect 375 137 376 138
rect 376 137 377 138
rect 377 137 378 138
rect 378 137 379 138
rect 379 137 380 138
rect 380 137 381 138
rect 381 137 382 138
rect 382 137 383 138
rect 383 137 384 138
rect 384 137 385 138
rect 385 137 386 138
rect 386 137 387 138
rect 387 137 388 138
rect 388 137 389 138
rect 389 137 390 138
rect 390 137 391 138
rect 391 137 392 138
rect 392 137 393 138
rect 393 137 394 138
rect 394 137 395 138
rect 395 137 396 138
rect 396 137 397 138
rect 397 137 398 138
rect 398 137 399 138
rect 399 137 400 138
rect 400 137 401 138
rect 401 137 402 138
rect 402 137 403 138
rect 403 137 404 138
rect 404 137 405 138
rect 405 137 406 138
rect 406 137 407 138
rect 407 137 408 138
rect 408 137 409 138
rect 409 137 410 138
rect 476 137 477 138
rect 477 137 478 138
rect 478 137 479 138
rect 479 137 480 138
rect 480 137 481 138
rect 481 137 482 138
rect 482 137 483 138
rect 483 137 484 138
rect 484 137 485 138
rect 485 137 486 138
rect 486 137 487 138
rect 487 137 488 138
rect 488 137 489 138
rect 489 137 490 138
rect 490 137 491 138
rect 491 137 492 138
rect 492 137 493 138
rect 493 137 494 138
rect 494 137 495 138
rect 495 137 496 138
rect 496 137 497 138
rect 497 137 498 138
rect 117 136 118 137
rect 118 136 119 137
rect 119 136 120 137
rect 120 136 121 137
rect 121 136 122 137
rect 122 136 123 137
rect 123 136 124 137
rect 124 136 125 137
rect 125 136 126 137
rect 126 136 127 137
rect 127 136 128 137
rect 128 136 129 137
rect 129 136 130 137
rect 130 136 131 137
rect 272 136 273 137
rect 273 136 274 137
rect 274 136 275 137
rect 275 136 276 137
rect 276 136 277 137
rect 277 136 278 137
rect 278 136 279 137
rect 300 136 301 137
rect 301 136 302 137
rect 302 136 303 137
rect 303 136 304 137
rect 304 136 305 137
rect 305 136 306 137
rect 306 136 307 137
rect 307 136 308 137
rect 308 136 309 137
rect 309 136 310 137
rect 310 136 311 137
rect 311 136 312 137
rect 312 136 313 137
rect 313 136 314 137
rect 336 136 337 137
rect 337 136 338 137
rect 338 136 339 137
rect 339 136 340 137
rect 340 136 341 137
rect 341 136 342 137
rect 342 136 343 137
rect 343 136 344 137
rect 344 136 345 137
rect 345 136 346 137
rect 346 136 347 137
rect 347 136 348 137
rect 362 136 363 137
rect 363 136 364 137
rect 364 136 365 137
rect 365 136 366 137
rect 366 136 367 137
rect 367 136 368 137
rect 368 136 369 137
rect 369 136 370 137
rect 370 136 371 137
rect 371 136 372 137
rect 372 136 373 137
rect 373 136 374 137
rect 374 136 375 137
rect 375 136 376 137
rect 376 136 377 137
rect 377 136 378 137
rect 378 136 379 137
rect 379 136 380 137
rect 380 136 381 137
rect 381 136 382 137
rect 382 136 383 137
rect 383 136 384 137
rect 384 136 385 137
rect 385 136 386 137
rect 386 136 387 137
rect 387 136 388 137
rect 388 136 389 137
rect 389 136 390 137
rect 390 136 391 137
rect 391 136 392 137
rect 392 136 393 137
rect 393 136 394 137
rect 394 136 395 137
rect 395 136 396 137
rect 396 136 397 137
rect 397 136 398 137
rect 398 136 399 137
rect 399 136 400 137
rect 400 136 401 137
rect 401 136 402 137
rect 402 136 403 137
rect 403 136 404 137
rect 404 136 405 137
rect 405 136 406 137
rect 406 136 407 137
rect 407 136 408 137
rect 408 136 409 137
rect 409 136 410 137
rect 474 136 475 137
rect 475 136 476 137
rect 476 136 477 137
rect 477 136 478 137
rect 478 136 479 137
rect 479 136 480 137
rect 480 136 481 137
rect 481 136 482 137
rect 482 136 483 137
rect 483 136 484 137
rect 484 136 485 137
rect 485 136 486 137
rect 486 136 487 137
rect 487 136 488 137
rect 488 136 489 137
rect 489 136 490 137
rect 490 136 491 137
rect 491 136 492 137
rect 492 136 493 137
rect 493 136 494 137
rect 494 136 495 137
rect 495 136 496 137
rect 496 136 497 137
rect 497 136 498 137
rect 118 135 119 136
rect 119 135 120 136
rect 120 135 121 136
rect 121 135 122 136
rect 122 135 123 136
rect 123 135 124 136
rect 124 135 125 136
rect 125 135 126 136
rect 126 135 127 136
rect 127 135 128 136
rect 128 135 129 136
rect 129 135 130 136
rect 130 135 131 136
rect 272 135 273 136
rect 273 135 274 136
rect 274 135 275 136
rect 275 135 276 136
rect 276 135 277 136
rect 302 135 303 136
rect 303 135 304 136
rect 304 135 305 136
rect 305 135 306 136
rect 306 135 307 136
rect 307 135 308 136
rect 308 135 309 136
rect 309 135 310 136
rect 310 135 311 136
rect 311 135 312 136
rect 312 135 313 136
rect 313 135 314 136
rect 336 135 337 136
rect 337 135 338 136
rect 338 135 339 136
rect 339 135 340 136
rect 340 135 341 136
rect 341 135 342 136
rect 342 135 343 136
rect 343 135 344 136
rect 344 135 345 136
rect 345 135 346 136
rect 362 135 363 136
rect 363 135 364 136
rect 364 135 365 136
rect 365 135 366 136
rect 366 135 367 136
rect 367 135 368 136
rect 368 135 369 136
rect 369 135 370 136
rect 370 135 371 136
rect 371 135 372 136
rect 372 135 373 136
rect 373 135 374 136
rect 374 135 375 136
rect 375 135 376 136
rect 376 135 377 136
rect 377 135 378 136
rect 378 135 379 136
rect 379 135 380 136
rect 380 135 381 136
rect 381 135 382 136
rect 382 135 383 136
rect 383 135 384 136
rect 384 135 385 136
rect 385 135 386 136
rect 386 135 387 136
rect 387 135 388 136
rect 388 135 389 136
rect 389 135 390 136
rect 390 135 391 136
rect 391 135 392 136
rect 392 135 393 136
rect 393 135 394 136
rect 394 135 395 136
rect 395 135 396 136
rect 396 135 397 136
rect 397 135 398 136
rect 398 135 399 136
rect 399 135 400 136
rect 400 135 401 136
rect 401 135 402 136
rect 402 135 403 136
rect 403 135 404 136
rect 404 135 405 136
rect 405 135 406 136
rect 406 135 407 136
rect 407 135 408 136
rect 408 135 409 136
rect 409 135 410 136
rect 474 135 475 136
rect 475 135 476 136
rect 476 135 477 136
rect 477 135 478 136
rect 478 135 479 136
rect 479 135 480 136
rect 480 135 481 136
rect 481 135 482 136
rect 482 135 483 136
rect 483 135 484 136
rect 484 135 485 136
rect 485 135 486 136
rect 486 135 487 136
rect 487 135 488 136
rect 488 135 489 136
rect 489 135 490 136
rect 490 135 491 136
rect 491 135 492 136
rect 492 135 493 136
rect 493 135 494 136
rect 494 135 495 136
rect 495 135 496 136
rect 118 134 119 135
rect 119 134 120 135
rect 120 134 121 135
rect 121 134 122 135
rect 122 134 123 135
rect 123 134 124 135
rect 124 134 125 135
rect 125 134 126 135
rect 126 134 127 135
rect 127 134 128 135
rect 128 134 129 135
rect 129 134 130 135
rect 130 134 131 135
rect 270 134 271 135
rect 271 134 272 135
rect 272 134 273 135
rect 273 134 274 135
rect 274 134 275 135
rect 275 134 276 135
rect 276 134 277 135
rect 302 134 303 135
rect 303 134 304 135
rect 304 134 305 135
rect 305 134 306 135
rect 306 134 307 135
rect 307 134 308 135
rect 308 134 309 135
rect 309 134 310 135
rect 310 134 311 135
rect 311 134 312 135
rect 312 134 313 135
rect 313 134 314 135
rect 336 134 337 135
rect 337 134 338 135
rect 338 134 339 135
rect 339 134 340 135
rect 340 134 341 135
rect 341 134 342 135
rect 342 134 343 135
rect 343 134 344 135
rect 344 134 345 135
rect 345 134 346 135
rect 360 134 361 135
rect 361 134 362 135
rect 362 134 363 135
rect 363 134 364 135
rect 364 134 365 135
rect 365 134 366 135
rect 366 134 367 135
rect 367 134 368 135
rect 368 134 369 135
rect 369 134 370 135
rect 370 134 371 135
rect 371 134 372 135
rect 372 134 373 135
rect 373 134 374 135
rect 374 134 375 135
rect 375 134 376 135
rect 376 134 377 135
rect 377 134 378 135
rect 378 134 379 135
rect 379 134 380 135
rect 380 134 381 135
rect 381 134 382 135
rect 382 134 383 135
rect 383 134 384 135
rect 384 134 385 135
rect 385 134 386 135
rect 386 134 387 135
rect 387 134 388 135
rect 388 134 389 135
rect 389 134 390 135
rect 390 134 391 135
rect 391 134 392 135
rect 392 134 393 135
rect 393 134 394 135
rect 394 134 395 135
rect 395 134 396 135
rect 396 134 397 135
rect 397 134 398 135
rect 398 134 399 135
rect 399 134 400 135
rect 400 134 401 135
rect 401 134 402 135
rect 402 134 403 135
rect 403 134 404 135
rect 404 134 405 135
rect 405 134 406 135
rect 406 134 407 135
rect 407 134 408 135
rect 408 134 409 135
rect 409 134 410 135
rect 472 134 473 135
rect 473 134 474 135
rect 474 134 475 135
rect 475 134 476 135
rect 476 134 477 135
rect 477 134 478 135
rect 478 134 479 135
rect 479 134 480 135
rect 480 134 481 135
rect 481 134 482 135
rect 482 134 483 135
rect 483 134 484 135
rect 484 134 485 135
rect 485 134 486 135
rect 486 134 487 135
rect 487 134 488 135
rect 488 134 489 135
rect 489 134 490 135
rect 490 134 491 135
rect 491 134 492 135
rect 492 134 493 135
rect 493 134 494 135
rect 494 134 495 135
rect 495 134 496 135
rect 118 133 119 134
rect 119 133 120 134
rect 120 133 121 134
rect 121 133 122 134
rect 122 133 123 134
rect 123 133 124 134
rect 124 133 125 134
rect 125 133 126 134
rect 126 133 127 134
rect 127 133 128 134
rect 128 133 129 134
rect 129 133 130 134
rect 130 133 131 134
rect 270 133 271 134
rect 271 133 272 134
rect 272 133 273 134
rect 273 133 274 134
rect 274 133 275 134
rect 275 133 276 134
rect 276 133 277 134
rect 302 133 303 134
rect 303 133 304 134
rect 304 133 305 134
rect 305 133 306 134
rect 306 133 307 134
rect 307 133 308 134
rect 308 133 309 134
rect 309 133 310 134
rect 310 133 311 134
rect 311 133 312 134
rect 312 133 313 134
rect 313 133 314 134
rect 336 133 337 134
rect 337 133 338 134
rect 338 133 339 134
rect 339 133 340 134
rect 340 133 341 134
rect 341 133 342 134
rect 342 133 343 134
rect 343 133 344 134
rect 344 133 345 134
rect 345 133 346 134
rect 360 133 361 134
rect 361 133 362 134
rect 362 133 363 134
rect 363 133 364 134
rect 364 133 365 134
rect 365 133 366 134
rect 366 133 367 134
rect 367 133 368 134
rect 368 133 369 134
rect 369 133 370 134
rect 370 133 371 134
rect 371 133 372 134
rect 372 133 373 134
rect 373 133 374 134
rect 374 133 375 134
rect 375 133 376 134
rect 376 133 377 134
rect 377 133 378 134
rect 378 133 379 134
rect 379 133 380 134
rect 380 133 381 134
rect 381 133 382 134
rect 382 133 383 134
rect 383 133 384 134
rect 384 133 385 134
rect 385 133 386 134
rect 386 133 387 134
rect 387 133 388 134
rect 388 133 389 134
rect 389 133 390 134
rect 390 133 391 134
rect 391 133 392 134
rect 392 133 393 134
rect 393 133 394 134
rect 394 133 395 134
rect 395 133 396 134
rect 396 133 397 134
rect 397 133 398 134
rect 398 133 399 134
rect 399 133 400 134
rect 400 133 401 134
rect 401 133 402 134
rect 402 133 403 134
rect 403 133 404 134
rect 404 133 405 134
rect 405 133 406 134
rect 406 133 407 134
rect 407 133 408 134
rect 408 133 409 134
rect 409 133 410 134
rect 472 133 473 134
rect 473 133 474 134
rect 474 133 475 134
rect 475 133 476 134
rect 476 133 477 134
rect 477 133 478 134
rect 478 133 479 134
rect 479 133 480 134
rect 480 133 481 134
rect 481 133 482 134
rect 482 133 483 134
rect 483 133 484 134
rect 484 133 485 134
rect 485 133 486 134
rect 486 133 487 134
rect 487 133 488 134
rect 488 133 489 134
rect 489 133 490 134
rect 490 133 491 134
rect 491 133 492 134
rect 118 132 119 133
rect 119 132 120 133
rect 120 132 121 133
rect 121 132 122 133
rect 122 132 123 133
rect 123 132 124 133
rect 124 132 125 133
rect 125 132 126 133
rect 126 132 127 133
rect 127 132 128 133
rect 128 132 129 133
rect 129 132 130 133
rect 130 132 131 133
rect 131 132 132 133
rect 132 132 133 133
rect 268 132 269 133
rect 269 132 270 133
rect 270 132 271 133
rect 271 132 272 133
rect 272 132 273 133
rect 273 132 274 133
rect 274 132 275 133
rect 275 132 276 133
rect 276 132 277 133
rect 302 132 303 133
rect 303 132 304 133
rect 304 132 305 133
rect 305 132 306 133
rect 306 132 307 133
rect 307 132 308 133
rect 308 132 309 133
rect 309 132 310 133
rect 310 132 311 133
rect 311 132 312 133
rect 312 132 313 133
rect 313 132 314 133
rect 314 132 315 133
rect 315 132 316 133
rect 336 132 337 133
rect 337 132 338 133
rect 338 132 339 133
rect 339 132 340 133
rect 340 132 341 133
rect 341 132 342 133
rect 342 132 343 133
rect 343 132 344 133
rect 344 132 345 133
rect 345 132 346 133
rect 358 132 359 133
rect 359 132 360 133
rect 360 132 361 133
rect 361 132 362 133
rect 362 132 363 133
rect 363 132 364 133
rect 364 132 365 133
rect 365 132 366 133
rect 366 132 367 133
rect 367 132 368 133
rect 368 132 369 133
rect 369 132 370 133
rect 370 132 371 133
rect 371 132 372 133
rect 372 132 373 133
rect 373 132 374 133
rect 374 132 375 133
rect 375 132 376 133
rect 376 132 377 133
rect 377 132 378 133
rect 378 132 379 133
rect 379 132 380 133
rect 380 132 381 133
rect 381 132 382 133
rect 382 132 383 133
rect 383 132 384 133
rect 384 132 385 133
rect 385 132 386 133
rect 386 132 387 133
rect 387 132 388 133
rect 388 132 389 133
rect 389 132 390 133
rect 390 132 391 133
rect 391 132 392 133
rect 392 132 393 133
rect 393 132 394 133
rect 394 132 395 133
rect 395 132 396 133
rect 396 132 397 133
rect 397 132 398 133
rect 398 132 399 133
rect 399 132 400 133
rect 400 132 401 133
rect 401 132 402 133
rect 402 132 403 133
rect 403 132 404 133
rect 404 132 405 133
rect 405 132 406 133
rect 406 132 407 133
rect 407 132 408 133
rect 408 132 409 133
rect 409 132 410 133
rect 471 132 472 133
rect 472 132 473 133
rect 473 132 474 133
rect 474 132 475 133
rect 475 132 476 133
rect 476 132 477 133
rect 477 132 478 133
rect 478 132 479 133
rect 479 132 480 133
rect 480 132 481 133
rect 481 132 482 133
rect 482 132 483 133
rect 483 132 484 133
rect 484 132 485 133
rect 485 132 486 133
rect 486 132 487 133
rect 487 132 488 133
rect 488 132 489 133
rect 489 132 490 133
rect 490 132 491 133
rect 491 132 492 133
rect 120 131 121 132
rect 121 131 122 132
rect 122 131 123 132
rect 123 131 124 132
rect 124 131 125 132
rect 125 131 126 132
rect 126 131 127 132
rect 127 131 128 132
rect 128 131 129 132
rect 129 131 130 132
rect 130 131 131 132
rect 131 131 132 132
rect 132 131 133 132
rect 268 131 269 132
rect 269 131 270 132
rect 270 131 271 132
rect 271 131 272 132
rect 272 131 273 132
rect 273 131 274 132
rect 274 131 275 132
rect 275 131 276 132
rect 276 131 277 132
rect 304 131 305 132
rect 305 131 306 132
rect 306 131 307 132
rect 307 131 308 132
rect 308 131 309 132
rect 309 131 310 132
rect 310 131 311 132
rect 311 131 312 132
rect 312 131 313 132
rect 313 131 314 132
rect 314 131 315 132
rect 315 131 316 132
rect 336 131 337 132
rect 337 131 338 132
rect 338 131 339 132
rect 339 131 340 132
rect 340 131 341 132
rect 341 131 342 132
rect 342 131 343 132
rect 343 131 344 132
rect 344 131 345 132
rect 345 131 346 132
rect 358 131 359 132
rect 359 131 360 132
rect 360 131 361 132
rect 361 131 362 132
rect 362 131 363 132
rect 363 131 364 132
rect 364 131 365 132
rect 365 131 366 132
rect 366 131 367 132
rect 367 131 368 132
rect 368 131 369 132
rect 369 131 370 132
rect 370 131 371 132
rect 371 131 372 132
rect 372 131 373 132
rect 373 131 374 132
rect 374 131 375 132
rect 375 131 376 132
rect 376 131 377 132
rect 377 131 378 132
rect 378 131 379 132
rect 379 131 380 132
rect 380 131 381 132
rect 381 131 382 132
rect 382 131 383 132
rect 383 131 384 132
rect 384 131 385 132
rect 385 131 386 132
rect 386 131 387 132
rect 387 131 388 132
rect 388 131 389 132
rect 389 131 390 132
rect 390 131 391 132
rect 391 131 392 132
rect 392 131 393 132
rect 393 131 394 132
rect 394 131 395 132
rect 395 131 396 132
rect 396 131 397 132
rect 397 131 398 132
rect 398 131 399 132
rect 399 131 400 132
rect 400 131 401 132
rect 401 131 402 132
rect 402 131 403 132
rect 403 131 404 132
rect 404 131 405 132
rect 405 131 406 132
rect 406 131 407 132
rect 407 131 408 132
rect 471 131 472 132
rect 472 131 473 132
rect 473 131 474 132
rect 474 131 475 132
rect 475 131 476 132
rect 476 131 477 132
rect 477 131 478 132
rect 478 131 479 132
rect 479 131 480 132
rect 480 131 481 132
rect 481 131 482 132
rect 482 131 483 132
rect 483 131 484 132
rect 484 131 485 132
rect 485 131 486 132
rect 486 131 487 132
rect 487 131 488 132
rect 488 131 489 132
rect 489 131 490 132
rect 490 131 491 132
rect 491 131 492 132
rect 120 130 121 131
rect 121 130 122 131
rect 122 130 123 131
rect 123 130 124 131
rect 124 130 125 131
rect 125 130 126 131
rect 126 130 127 131
rect 127 130 128 131
rect 128 130 129 131
rect 129 130 130 131
rect 130 130 131 131
rect 131 130 132 131
rect 132 130 133 131
rect 133 130 134 131
rect 268 130 269 131
rect 269 130 270 131
rect 270 130 271 131
rect 271 130 272 131
rect 272 130 273 131
rect 273 130 274 131
rect 274 130 275 131
rect 275 130 276 131
rect 276 130 277 131
rect 302 130 303 131
rect 303 130 304 131
rect 304 130 305 131
rect 305 130 306 131
rect 306 130 307 131
rect 307 130 308 131
rect 308 130 309 131
rect 309 130 310 131
rect 310 130 311 131
rect 311 130 312 131
rect 312 130 313 131
rect 313 130 314 131
rect 314 130 315 131
rect 315 130 316 131
rect 336 130 337 131
rect 337 130 338 131
rect 338 130 339 131
rect 339 130 340 131
rect 340 130 341 131
rect 341 130 342 131
rect 342 130 343 131
rect 343 130 344 131
rect 344 130 345 131
rect 345 130 346 131
rect 358 130 359 131
rect 359 130 360 131
rect 360 130 361 131
rect 361 130 362 131
rect 362 130 363 131
rect 363 130 364 131
rect 364 130 365 131
rect 365 130 366 131
rect 366 130 367 131
rect 367 130 368 131
rect 368 130 369 131
rect 369 130 370 131
rect 370 130 371 131
rect 371 130 372 131
rect 372 130 373 131
rect 373 130 374 131
rect 374 130 375 131
rect 375 130 376 131
rect 376 130 377 131
rect 377 130 378 131
rect 378 130 379 131
rect 379 130 380 131
rect 380 130 381 131
rect 381 130 382 131
rect 382 130 383 131
rect 383 130 384 131
rect 384 130 385 131
rect 385 130 386 131
rect 386 130 387 131
rect 387 130 388 131
rect 388 130 389 131
rect 389 130 390 131
rect 390 130 391 131
rect 391 130 392 131
rect 392 130 393 131
rect 393 130 394 131
rect 394 130 395 131
rect 395 130 396 131
rect 396 130 397 131
rect 397 130 398 131
rect 398 130 399 131
rect 399 130 400 131
rect 400 130 401 131
rect 401 130 402 131
rect 402 130 403 131
rect 403 130 404 131
rect 404 130 405 131
rect 405 130 406 131
rect 406 130 407 131
rect 407 130 408 131
rect 469 130 470 131
rect 470 130 471 131
rect 471 130 472 131
rect 472 130 473 131
rect 473 130 474 131
rect 474 130 475 131
rect 475 130 476 131
rect 476 130 477 131
rect 477 130 478 131
rect 478 130 479 131
rect 479 130 480 131
rect 480 130 481 131
rect 481 130 482 131
rect 482 130 483 131
rect 483 130 484 131
rect 484 130 485 131
rect 485 130 486 131
rect 486 130 487 131
rect 487 130 488 131
rect 488 130 489 131
rect 489 130 490 131
rect 490 130 491 131
rect 491 130 492 131
rect 120 129 121 130
rect 121 129 122 130
rect 122 129 123 130
rect 123 129 124 130
rect 124 129 125 130
rect 125 129 126 130
rect 126 129 127 130
rect 127 129 128 130
rect 128 129 129 130
rect 129 129 130 130
rect 130 129 131 130
rect 131 129 132 130
rect 132 129 133 130
rect 133 129 134 130
rect 268 129 269 130
rect 269 129 270 130
rect 270 129 271 130
rect 271 129 272 130
rect 272 129 273 130
rect 273 129 274 130
rect 274 129 275 130
rect 302 129 303 130
rect 303 129 304 130
rect 304 129 305 130
rect 305 129 306 130
rect 306 129 307 130
rect 307 129 308 130
rect 308 129 309 130
rect 309 129 310 130
rect 310 129 311 130
rect 311 129 312 130
rect 312 129 313 130
rect 313 129 314 130
rect 314 129 315 130
rect 315 129 316 130
rect 336 129 337 130
rect 337 129 338 130
rect 338 129 339 130
rect 339 129 340 130
rect 340 129 341 130
rect 341 129 342 130
rect 342 129 343 130
rect 343 129 344 130
rect 344 129 345 130
rect 345 129 346 130
rect 469 129 470 130
rect 470 129 471 130
rect 471 129 472 130
rect 472 129 473 130
rect 473 129 474 130
rect 474 129 475 130
rect 475 129 476 130
rect 476 129 477 130
rect 477 129 478 130
rect 478 129 479 130
rect 479 129 480 130
rect 480 129 481 130
rect 481 129 482 130
rect 482 129 483 130
rect 483 129 484 130
rect 484 129 485 130
rect 485 129 486 130
rect 486 129 487 130
rect 487 129 488 130
rect 488 129 489 130
rect 489 129 490 130
rect 120 128 121 129
rect 121 128 122 129
rect 122 128 123 129
rect 123 128 124 129
rect 124 128 125 129
rect 125 128 126 129
rect 126 128 127 129
rect 127 128 128 129
rect 128 128 129 129
rect 129 128 130 129
rect 130 128 131 129
rect 131 128 132 129
rect 132 128 133 129
rect 133 128 134 129
rect 268 128 269 129
rect 269 128 270 129
rect 270 128 271 129
rect 271 128 272 129
rect 272 128 273 129
rect 273 128 274 129
rect 274 128 275 129
rect 302 128 303 129
rect 303 128 304 129
rect 304 128 305 129
rect 305 128 306 129
rect 306 128 307 129
rect 307 128 308 129
rect 308 128 309 129
rect 309 128 310 129
rect 310 128 311 129
rect 311 128 312 129
rect 312 128 313 129
rect 313 128 314 129
rect 314 128 315 129
rect 315 128 316 129
rect 336 128 337 129
rect 337 128 338 129
rect 338 128 339 129
rect 339 128 340 129
rect 340 128 341 129
rect 341 128 342 129
rect 342 128 343 129
rect 343 128 344 129
rect 344 128 345 129
rect 345 128 346 129
rect 469 128 470 129
rect 470 128 471 129
rect 471 128 472 129
rect 472 128 473 129
rect 473 128 474 129
rect 474 128 475 129
rect 475 128 476 129
rect 476 128 477 129
rect 477 128 478 129
rect 478 128 479 129
rect 479 128 480 129
rect 480 128 481 129
rect 481 128 482 129
rect 482 128 483 129
rect 483 128 484 129
rect 484 128 485 129
rect 485 128 486 129
rect 486 128 487 129
rect 487 128 488 129
rect 488 128 489 129
rect 489 128 490 129
rect 120 127 121 128
rect 121 127 122 128
rect 122 127 123 128
rect 123 127 124 128
rect 124 127 125 128
rect 125 127 126 128
rect 126 127 127 128
rect 127 127 128 128
rect 128 127 129 128
rect 129 127 130 128
rect 130 127 131 128
rect 131 127 132 128
rect 132 127 133 128
rect 133 127 134 128
rect 265 127 266 128
rect 266 127 267 128
rect 267 127 268 128
rect 268 127 269 128
rect 269 127 270 128
rect 270 127 271 128
rect 271 127 272 128
rect 272 127 273 128
rect 273 127 274 128
rect 274 127 275 128
rect 275 127 276 128
rect 276 127 277 128
rect 302 127 303 128
rect 303 127 304 128
rect 304 127 305 128
rect 305 127 306 128
rect 306 127 307 128
rect 307 127 308 128
rect 308 127 309 128
rect 309 127 310 128
rect 310 127 311 128
rect 311 127 312 128
rect 312 127 313 128
rect 313 127 314 128
rect 314 127 315 128
rect 315 127 316 128
rect 316 127 317 128
rect 317 127 318 128
rect 318 127 319 128
rect 319 127 320 128
rect 336 127 337 128
rect 337 127 338 128
rect 338 127 339 128
rect 339 127 340 128
rect 340 127 341 128
rect 341 127 342 128
rect 342 127 343 128
rect 343 127 344 128
rect 344 127 345 128
rect 345 127 346 128
rect 346 127 347 128
rect 347 127 348 128
rect 465 127 466 128
rect 466 127 467 128
rect 467 127 468 128
rect 468 127 469 128
rect 469 127 470 128
rect 470 127 471 128
rect 471 127 472 128
rect 472 127 473 128
rect 473 127 474 128
rect 474 127 475 128
rect 475 127 476 128
rect 476 127 477 128
rect 477 127 478 128
rect 478 127 479 128
rect 479 127 480 128
rect 480 127 481 128
rect 481 127 482 128
rect 482 127 483 128
rect 483 127 484 128
rect 484 127 485 128
rect 485 127 486 128
rect 486 127 487 128
rect 487 127 488 128
rect 488 127 489 128
rect 489 127 490 128
rect 122 126 123 127
rect 123 126 124 127
rect 124 126 125 127
rect 125 126 126 127
rect 126 126 127 127
rect 127 126 128 127
rect 128 126 129 127
rect 129 126 130 127
rect 130 126 131 127
rect 131 126 132 127
rect 132 126 133 127
rect 133 126 134 127
rect 265 126 266 127
rect 266 126 267 127
rect 267 126 268 127
rect 268 126 269 127
rect 269 126 270 127
rect 270 126 271 127
rect 271 126 272 127
rect 272 126 273 127
rect 273 126 274 127
rect 274 126 275 127
rect 275 126 276 127
rect 276 126 277 127
rect 302 126 303 127
rect 303 126 304 127
rect 304 126 305 127
rect 305 126 306 127
rect 306 126 307 127
rect 307 126 308 127
rect 308 126 309 127
rect 309 126 310 127
rect 310 126 311 127
rect 311 126 312 127
rect 312 126 313 127
rect 313 126 314 127
rect 314 126 315 127
rect 315 126 316 127
rect 316 126 317 127
rect 317 126 318 127
rect 318 126 319 127
rect 319 126 320 127
rect 336 126 337 127
rect 337 126 338 127
rect 338 126 339 127
rect 339 126 340 127
rect 340 126 341 127
rect 341 126 342 127
rect 342 126 343 127
rect 343 126 344 127
rect 344 126 345 127
rect 345 126 346 127
rect 346 126 347 127
rect 347 126 348 127
rect 465 126 466 127
rect 466 126 467 127
rect 467 126 468 127
rect 468 126 469 127
rect 469 126 470 127
rect 470 126 471 127
rect 471 126 472 127
rect 472 126 473 127
rect 473 126 474 127
rect 474 126 475 127
rect 475 126 476 127
rect 476 126 477 127
rect 477 126 478 127
rect 478 126 479 127
rect 479 126 480 127
rect 480 126 481 127
rect 481 126 482 127
rect 482 126 483 127
rect 483 126 484 127
rect 484 126 485 127
rect 485 126 486 127
rect 486 126 487 127
rect 487 126 488 127
rect 122 125 123 126
rect 123 125 124 126
rect 124 125 125 126
rect 125 125 126 126
rect 126 125 127 126
rect 127 125 128 126
rect 128 125 129 126
rect 129 125 130 126
rect 130 125 131 126
rect 131 125 132 126
rect 132 125 133 126
rect 133 125 134 126
rect 134 125 135 126
rect 135 125 136 126
rect 261 125 262 126
rect 262 125 263 126
rect 263 125 264 126
rect 264 125 265 126
rect 265 125 266 126
rect 266 125 267 126
rect 267 125 268 126
rect 268 125 269 126
rect 269 125 270 126
rect 270 125 271 126
rect 271 125 272 126
rect 272 125 273 126
rect 273 125 274 126
rect 274 125 275 126
rect 275 125 276 126
rect 276 125 277 126
rect 277 125 278 126
rect 278 125 279 126
rect 279 125 280 126
rect 280 125 281 126
rect 281 125 282 126
rect 296 125 297 126
rect 297 125 298 126
rect 298 125 299 126
rect 299 125 300 126
rect 300 125 301 126
rect 301 125 302 126
rect 302 125 303 126
rect 303 125 304 126
rect 304 125 305 126
rect 305 125 306 126
rect 306 125 307 126
rect 307 125 308 126
rect 308 125 309 126
rect 309 125 310 126
rect 310 125 311 126
rect 311 125 312 126
rect 312 125 313 126
rect 313 125 314 126
rect 314 125 315 126
rect 315 125 316 126
rect 316 125 317 126
rect 317 125 318 126
rect 318 125 319 126
rect 319 125 320 126
rect 320 125 321 126
rect 321 125 322 126
rect 322 125 323 126
rect 323 125 324 126
rect 336 125 337 126
rect 337 125 338 126
rect 338 125 339 126
rect 339 125 340 126
rect 340 125 341 126
rect 341 125 342 126
rect 342 125 343 126
rect 343 125 344 126
rect 344 125 345 126
rect 345 125 346 126
rect 346 125 347 126
rect 347 125 348 126
rect 463 125 464 126
rect 464 125 465 126
rect 465 125 466 126
rect 466 125 467 126
rect 467 125 468 126
rect 468 125 469 126
rect 469 125 470 126
rect 470 125 471 126
rect 471 125 472 126
rect 472 125 473 126
rect 473 125 474 126
rect 474 125 475 126
rect 475 125 476 126
rect 476 125 477 126
rect 477 125 478 126
rect 478 125 479 126
rect 479 125 480 126
rect 480 125 481 126
rect 481 125 482 126
rect 482 125 483 126
rect 483 125 484 126
rect 484 125 485 126
rect 485 125 486 126
rect 486 125 487 126
rect 487 125 488 126
rect 124 124 125 125
rect 125 124 126 125
rect 126 124 127 125
rect 127 124 128 125
rect 128 124 129 125
rect 129 124 130 125
rect 130 124 131 125
rect 131 124 132 125
rect 132 124 133 125
rect 133 124 134 125
rect 134 124 135 125
rect 135 124 136 125
rect 261 124 262 125
rect 262 124 263 125
rect 263 124 264 125
rect 264 124 265 125
rect 265 124 266 125
rect 266 124 267 125
rect 267 124 268 125
rect 268 124 269 125
rect 269 124 270 125
rect 270 124 271 125
rect 271 124 272 125
rect 272 124 273 125
rect 273 124 274 125
rect 274 124 275 125
rect 275 124 276 125
rect 276 124 277 125
rect 277 124 278 125
rect 278 124 279 125
rect 279 124 280 125
rect 280 124 281 125
rect 281 124 282 125
rect 296 124 297 125
rect 297 124 298 125
rect 298 124 299 125
rect 299 124 300 125
rect 300 124 301 125
rect 301 124 302 125
rect 302 124 303 125
rect 303 124 304 125
rect 304 124 305 125
rect 305 124 306 125
rect 306 124 307 125
rect 307 124 308 125
rect 308 124 309 125
rect 309 124 310 125
rect 310 124 311 125
rect 311 124 312 125
rect 312 124 313 125
rect 313 124 314 125
rect 314 124 315 125
rect 315 124 316 125
rect 316 124 317 125
rect 317 124 318 125
rect 318 124 319 125
rect 319 124 320 125
rect 320 124 321 125
rect 321 124 322 125
rect 322 124 323 125
rect 323 124 324 125
rect 336 124 337 125
rect 337 124 338 125
rect 338 124 339 125
rect 339 124 340 125
rect 340 124 341 125
rect 341 124 342 125
rect 342 124 343 125
rect 343 124 344 125
rect 344 124 345 125
rect 345 124 346 125
rect 346 124 347 125
rect 347 124 348 125
rect 463 124 464 125
rect 464 124 465 125
rect 465 124 466 125
rect 466 124 467 125
rect 467 124 468 125
rect 468 124 469 125
rect 469 124 470 125
rect 470 124 471 125
rect 471 124 472 125
rect 472 124 473 125
rect 473 124 474 125
rect 474 124 475 125
rect 475 124 476 125
rect 476 124 477 125
rect 477 124 478 125
rect 478 124 479 125
rect 479 124 480 125
rect 480 124 481 125
rect 481 124 482 125
rect 482 124 483 125
rect 483 124 484 125
rect 484 124 485 125
rect 485 124 486 125
rect 486 124 487 125
rect 124 123 125 124
rect 125 123 126 124
rect 126 123 127 124
rect 127 123 128 124
rect 128 123 129 124
rect 129 123 130 124
rect 130 123 131 124
rect 131 123 132 124
rect 132 123 133 124
rect 133 123 134 124
rect 134 123 135 124
rect 135 123 136 124
rect 136 123 137 124
rect 137 123 138 124
rect 261 123 262 124
rect 262 123 263 124
rect 263 123 264 124
rect 264 123 265 124
rect 265 123 266 124
rect 266 123 267 124
rect 267 123 268 124
rect 268 123 269 124
rect 269 123 270 124
rect 270 123 271 124
rect 271 123 272 124
rect 272 123 273 124
rect 273 123 274 124
rect 274 123 275 124
rect 275 123 276 124
rect 276 123 277 124
rect 277 123 278 124
rect 278 123 279 124
rect 279 123 280 124
rect 280 123 281 124
rect 281 123 282 124
rect 296 123 297 124
rect 297 123 298 124
rect 298 123 299 124
rect 299 123 300 124
rect 300 123 301 124
rect 301 123 302 124
rect 302 123 303 124
rect 303 123 304 124
rect 304 123 305 124
rect 305 123 306 124
rect 306 123 307 124
rect 307 123 308 124
rect 308 123 309 124
rect 309 123 310 124
rect 310 123 311 124
rect 311 123 312 124
rect 312 123 313 124
rect 313 123 314 124
rect 314 123 315 124
rect 315 123 316 124
rect 316 123 317 124
rect 317 123 318 124
rect 318 123 319 124
rect 319 123 320 124
rect 320 123 321 124
rect 321 123 322 124
rect 322 123 323 124
rect 323 123 324 124
rect 336 123 337 124
rect 337 123 338 124
rect 338 123 339 124
rect 339 123 340 124
rect 340 123 341 124
rect 341 123 342 124
rect 342 123 343 124
rect 343 123 344 124
rect 344 123 345 124
rect 345 123 346 124
rect 346 123 347 124
rect 347 123 348 124
rect 459 123 460 124
rect 460 123 461 124
rect 461 123 462 124
rect 462 123 463 124
rect 463 123 464 124
rect 464 123 465 124
rect 465 123 466 124
rect 466 123 467 124
rect 467 123 468 124
rect 468 123 469 124
rect 469 123 470 124
rect 470 123 471 124
rect 471 123 472 124
rect 472 123 473 124
rect 473 123 474 124
rect 474 123 475 124
rect 475 123 476 124
rect 476 123 477 124
rect 477 123 478 124
rect 478 123 479 124
rect 479 123 480 124
rect 480 123 481 124
rect 481 123 482 124
rect 482 123 483 124
rect 483 123 484 124
rect 484 123 485 124
rect 485 123 486 124
rect 486 123 487 124
rect 124 122 125 123
rect 125 122 126 123
rect 126 122 127 123
rect 127 122 128 123
rect 128 122 129 123
rect 129 122 130 123
rect 130 122 131 123
rect 131 122 132 123
rect 132 122 133 123
rect 133 122 134 123
rect 134 122 135 123
rect 135 122 136 123
rect 136 122 137 123
rect 137 122 138 123
rect 265 122 266 123
rect 266 122 267 123
rect 270 122 271 123
rect 271 122 272 123
rect 272 122 273 123
rect 276 122 277 123
rect 277 122 278 123
rect 278 122 279 123
rect 300 122 301 123
rect 301 122 302 123
rect 302 122 303 123
rect 304 122 305 123
rect 305 122 306 123
rect 306 122 307 123
rect 311 122 312 123
rect 312 122 313 123
rect 313 122 314 123
rect 314 122 315 123
rect 315 122 316 123
rect 336 122 337 123
rect 337 122 338 123
rect 338 122 339 123
rect 339 122 340 123
rect 340 122 341 123
rect 341 122 342 123
rect 342 122 343 123
rect 343 122 344 123
rect 344 122 345 123
rect 345 122 346 123
rect 459 122 460 123
rect 460 122 461 123
rect 461 122 462 123
rect 462 122 463 123
rect 463 122 464 123
rect 464 122 465 123
rect 465 122 466 123
rect 466 122 467 123
rect 467 122 468 123
rect 468 122 469 123
rect 469 122 470 123
rect 470 122 471 123
rect 471 122 472 123
rect 472 122 473 123
rect 473 122 474 123
rect 474 122 475 123
rect 475 122 476 123
rect 476 122 477 123
rect 477 122 478 123
rect 478 122 479 123
rect 479 122 480 123
rect 480 122 481 123
rect 481 122 482 123
rect 482 122 483 123
rect 124 121 125 122
rect 125 121 126 122
rect 126 121 127 122
rect 127 121 128 122
rect 128 121 129 122
rect 129 121 130 122
rect 130 121 131 122
rect 131 121 132 122
rect 132 121 133 122
rect 133 121 134 122
rect 134 121 135 122
rect 135 121 136 122
rect 136 121 137 122
rect 137 121 138 122
rect 138 121 139 122
rect 139 121 140 122
rect 265 121 266 122
rect 266 121 267 122
rect 270 121 271 122
rect 271 121 272 122
rect 272 121 273 122
rect 276 121 277 122
rect 277 121 278 122
rect 278 121 279 122
rect 300 121 301 122
rect 301 121 302 122
rect 302 121 303 122
rect 304 121 305 122
rect 305 121 306 122
rect 306 121 307 122
rect 311 121 312 122
rect 312 121 313 122
rect 313 121 314 122
rect 314 121 315 122
rect 315 121 316 122
rect 336 121 337 122
rect 337 121 338 122
rect 338 121 339 122
rect 339 121 340 122
rect 340 121 341 122
rect 341 121 342 122
rect 342 121 343 122
rect 343 121 344 122
rect 344 121 345 122
rect 345 121 346 122
rect 457 121 458 122
rect 458 121 459 122
rect 459 121 460 122
rect 460 121 461 122
rect 461 121 462 122
rect 462 121 463 122
rect 463 121 464 122
rect 464 121 465 122
rect 465 121 466 122
rect 466 121 467 122
rect 467 121 468 122
rect 468 121 469 122
rect 469 121 470 122
rect 470 121 471 122
rect 471 121 472 122
rect 472 121 473 122
rect 473 121 474 122
rect 474 121 475 122
rect 475 121 476 122
rect 476 121 477 122
rect 477 121 478 122
rect 478 121 479 122
rect 479 121 480 122
rect 480 121 481 122
rect 481 121 482 122
rect 482 121 483 122
rect 126 120 127 121
rect 127 120 128 121
rect 128 120 129 121
rect 129 120 130 121
rect 130 120 131 121
rect 131 120 132 121
rect 132 120 133 121
rect 133 120 134 121
rect 134 120 135 121
rect 135 120 136 121
rect 136 120 137 121
rect 137 120 138 121
rect 138 120 139 121
rect 139 120 140 121
rect 336 120 337 121
rect 337 120 338 121
rect 338 120 339 121
rect 339 120 340 121
rect 340 120 341 121
rect 341 120 342 121
rect 342 120 343 121
rect 343 120 344 121
rect 344 120 345 121
rect 345 120 346 121
rect 457 120 458 121
rect 458 120 459 121
rect 459 120 460 121
rect 460 120 461 121
rect 461 120 462 121
rect 462 120 463 121
rect 463 120 464 121
rect 464 120 465 121
rect 465 120 466 121
rect 466 120 467 121
rect 467 120 468 121
rect 468 120 469 121
rect 469 120 470 121
rect 470 120 471 121
rect 471 120 472 121
rect 472 120 473 121
rect 473 120 474 121
rect 474 120 475 121
rect 475 120 476 121
rect 476 120 477 121
rect 477 120 478 121
rect 478 120 479 121
rect 479 120 480 121
rect 480 120 481 121
rect 126 119 127 120
rect 127 119 128 120
rect 128 119 129 120
rect 129 119 130 120
rect 130 119 131 120
rect 131 119 132 120
rect 132 119 133 120
rect 133 119 134 120
rect 134 119 135 120
rect 135 119 136 120
rect 136 119 137 120
rect 137 119 138 120
rect 138 119 139 120
rect 139 119 140 120
rect 336 119 337 120
rect 337 119 338 120
rect 338 119 339 120
rect 339 119 340 120
rect 340 119 341 120
rect 341 119 342 120
rect 342 119 343 120
rect 343 119 344 120
rect 344 119 345 120
rect 345 119 346 120
rect 346 119 347 120
rect 347 119 348 120
rect 456 119 457 120
rect 457 119 458 120
rect 458 119 459 120
rect 459 119 460 120
rect 460 119 461 120
rect 461 119 462 120
rect 462 119 463 120
rect 463 119 464 120
rect 464 119 465 120
rect 465 119 466 120
rect 466 119 467 120
rect 467 119 468 120
rect 468 119 469 120
rect 469 119 470 120
rect 470 119 471 120
rect 471 119 472 120
rect 472 119 473 120
rect 473 119 474 120
rect 474 119 475 120
rect 475 119 476 120
rect 476 119 477 120
rect 477 119 478 120
rect 478 119 479 120
rect 479 119 480 120
rect 480 119 481 120
rect 128 118 129 119
rect 129 118 130 119
rect 130 118 131 119
rect 131 118 132 119
rect 132 118 133 119
rect 133 118 134 119
rect 134 118 135 119
rect 135 118 136 119
rect 136 118 137 119
rect 137 118 138 119
rect 138 118 139 119
rect 139 118 140 119
rect 336 118 337 119
rect 337 118 338 119
rect 338 118 339 119
rect 339 118 340 119
rect 340 118 341 119
rect 341 118 342 119
rect 342 118 343 119
rect 343 118 344 119
rect 344 118 345 119
rect 345 118 346 119
rect 346 118 347 119
rect 347 118 348 119
rect 456 118 457 119
rect 457 118 458 119
rect 458 118 459 119
rect 459 118 460 119
rect 460 118 461 119
rect 461 118 462 119
rect 462 118 463 119
rect 463 118 464 119
rect 464 118 465 119
rect 465 118 466 119
rect 466 118 467 119
rect 467 118 468 119
rect 468 118 469 119
rect 469 118 470 119
rect 470 118 471 119
rect 471 118 472 119
rect 472 118 473 119
rect 473 118 474 119
rect 474 118 475 119
rect 475 118 476 119
rect 476 118 477 119
rect 477 118 478 119
rect 478 118 479 119
rect 128 117 129 118
rect 129 117 130 118
rect 130 117 131 118
rect 131 117 132 118
rect 132 117 133 118
rect 133 117 134 118
rect 134 117 135 118
rect 135 117 136 118
rect 136 117 137 118
rect 137 117 138 118
rect 138 117 139 118
rect 139 117 140 118
rect 140 117 141 118
rect 141 117 142 118
rect 336 117 337 118
rect 337 117 338 118
rect 338 117 339 118
rect 339 117 340 118
rect 340 117 341 118
rect 341 117 342 118
rect 342 117 343 118
rect 343 117 344 118
rect 344 117 345 118
rect 345 117 346 118
rect 346 117 347 118
rect 347 117 348 118
rect 454 117 455 118
rect 455 117 456 118
rect 456 117 457 118
rect 457 117 458 118
rect 458 117 459 118
rect 459 117 460 118
rect 460 117 461 118
rect 461 117 462 118
rect 462 117 463 118
rect 463 117 464 118
rect 464 117 465 118
rect 465 117 466 118
rect 466 117 467 118
rect 467 117 468 118
rect 468 117 469 118
rect 469 117 470 118
rect 470 117 471 118
rect 471 117 472 118
rect 472 117 473 118
rect 473 117 474 118
rect 474 117 475 118
rect 475 117 476 118
rect 476 117 477 118
rect 477 117 478 118
rect 478 117 479 118
rect 128 116 129 117
rect 129 116 130 117
rect 130 116 131 117
rect 131 116 132 117
rect 132 116 133 117
rect 133 116 134 117
rect 134 116 135 117
rect 135 116 136 117
rect 136 116 137 117
rect 137 116 138 117
rect 138 116 139 117
rect 139 116 140 117
rect 140 116 141 117
rect 141 116 142 117
rect 336 116 337 117
rect 337 116 338 117
rect 338 116 339 117
rect 339 116 340 117
rect 340 116 341 117
rect 341 116 342 117
rect 342 116 343 117
rect 343 116 344 117
rect 344 116 345 117
rect 345 116 346 117
rect 454 116 455 117
rect 455 116 456 117
rect 456 116 457 117
rect 457 116 458 117
rect 458 116 459 117
rect 459 116 460 117
rect 460 116 461 117
rect 461 116 462 117
rect 462 116 463 117
rect 463 116 464 117
rect 464 116 465 117
rect 465 116 466 117
rect 466 116 467 117
rect 467 116 468 117
rect 468 116 469 117
rect 469 116 470 117
rect 470 116 471 117
rect 471 116 472 117
rect 472 116 473 117
rect 473 116 474 117
rect 474 116 475 117
rect 475 116 476 117
rect 476 116 477 117
rect 128 115 129 116
rect 129 115 130 116
rect 130 115 131 116
rect 131 115 132 116
rect 132 115 133 116
rect 133 115 134 116
rect 134 115 135 116
rect 135 115 136 116
rect 136 115 137 116
rect 137 115 138 116
rect 138 115 139 116
rect 139 115 140 116
rect 140 115 141 116
rect 141 115 142 116
rect 142 115 143 116
rect 143 115 144 116
rect 336 115 337 116
rect 337 115 338 116
rect 338 115 339 116
rect 339 115 340 116
rect 340 115 341 116
rect 341 115 342 116
rect 342 115 343 116
rect 343 115 344 116
rect 344 115 345 116
rect 345 115 346 116
rect 346 115 347 116
rect 347 115 348 116
rect 450 115 451 116
rect 451 115 452 116
rect 452 115 453 116
rect 453 115 454 116
rect 454 115 455 116
rect 455 115 456 116
rect 456 115 457 116
rect 457 115 458 116
rect 458 115 459 116
rect 459 115 460 116
rect 460 115 461 116
rect 461 115 462 116
rect 462 115 463 116
rect 463 115 464 116
rect 464 115 465 116
rect 465 115 466 116
rect 466 115 467 116
rect 467 115 468 116
rect 468 115 469 116
rect 469 115 470 116
rect 470 115 471 116
rect 471 115 472 116
rect 472 115 473 116
rect 473 115 474 116
rect 474 115 475 116
rect 475 115 476 116
rect 476 115 477 116
rect 130 114 131 115
rect 131 114 132 115
rect 132 114 133 115
rect 133 114 134 115
rect 134 114 135 115
rect 135 114 136 115
rect 136 114 137 115
rect 137 114 138 115
rect 138 114 139 115
rect 139 114 140 115
rect 140 114 141 115
rect 141 114 142 115
rect 142 114 143 115
rect 143 114 144 115
rect 336 114 337 115
rect 337 114 338 115
rect 338 114 339 115
rect 339 114 340 115
rect 340 114 341 115
rect 341 114 342 115
rect 342 114 343 115
rect 343 114 344 115
rect 344 114 345 115
rect 345 114 346 115
rect 346 114 347 115
rect 347 114 348 115
rect 450 114 451 115
rect 451 114 452 115
rect 452 114 453 115
rect 453 114 454 115
rect 454 114 455 115
rect 455 114 456 115
rect 456 114 457 115
rect 457 114 458 115
rect 458 114 459 115
rect 459 114 460 115
rect 460 114 461 115
rect 461 114 462 115
rect 462 114 463 115
rect 463 114 464 115
rect 464 114 465 115
rect 465 114 466 115
rect 466 114 467 115
rect 467 114 468 115
rect 468 114 469 115
rect 469 114 470 115
rect 470 114 471 115
rect 471 114 472 115
rect 472 114 473 115
rect 473 114 474 115
rect 474 114 475 115
rect 130 113 131 114
rect 131 113 132 114
rect 132 113 133 114
rect 133 113 134 114
rect 134 113 135 114
rect 135 113 136 114
rect 136 113 137 114
rect 137 113 138 114
rect 138 113 139 114
rect 139 113 140 114
rect 140 113 141 114
rect 141 113 142 114
rect 142 113 143 114
rect 143 113 144 114
rect 144 113 145 114
rect 145 113 146 114
rect 332 113 333 114
rect 333 113 334 114
rect 334 113 335 114
rect 335 113 336 114
rect 336 113 337 114
rect 337 113 338 114
rect 338 113 339 114
rect 339 113 340 114
rect 340 113 341 114
rect 341 113 342 114
rect 342 113 343 114
rect 343 113 344 114
rect 344 113 345 114
rect 345 113 346 114
rect 346 113 347 114
rect 347 113 348 114
rect 348 113 349 114
rect 349 113 350 114
rect 448 113 449 114
rect 449 113 450 114
rect 450 113 451 114
rect 451 113 452 114
rect 452 113 453 114
rect 453 113 454 114
rect 454 113 455 114
rect 455 113 456 114
rect 456 113 457 114
rect 457 113 458 114
rect 458 113 459 114
rect 459 113 460 114
rect 460 113 461 114
rect 461 113 462 114
rect 462 113 463 114
rect 463 113 464 114
rect 464 113 465 114
rect 465 113 466 114
rect 466 113 467 114
rect 467 113 468 114
rect 468 113 469 114
rect 469 113 470 114
rect 470 113 471 114
rect 471 113 472 114
rect 472 113 473 114
rect 473 113 474 114
rect 474 113 475 114
rect 132 112 133 113
rect 133 112 134 113
rect 134 112 135 113
rect 135 112 136 113
rect 136 112 137 113
rect 137 112 138 113
rect 138 112 139 113
rect 139 112 140 113
rect 140 112 141 113
rect 141 112 142 113
rect 142 112 143 113
rect 143 112 144 113
rect 144 112 145 113
rect 145 112 146 113
rect 332 112 333 113
rect 333 112 334 113
rect 334 112 335 113
rect 335 112 336 113
rect 336 112 337 113
rect 337 112 338 113
rect 338 112 339 113
rect 339 112 340 113
rect 340 112 341 113
rect 341 112 342 113
rect 342 112 343 113
rect 343 112 344 113
rect 344 112 345 113
rect 345 112 346 113
rect 346 112 347 113
rect 347 112 348 113
rect 348 112 349 113
rect 349 112 350 113
rect 448 112 449 113
rect 449 112 450 113
rect 450 112 451 113
rect 451 112 452 113
rect 452 112 453 113
rect 453 112 454 113
rect 454 112 455 113
rect 455 112 456 113
rect 456 112 457 113
rect 457 112 458 113
rect 458 112 459 113
rect 459 112 460 113
rect 460 112 461 113
rect 461 112 462 113
rect 462 112 463 113
rect 463 112 464 113
rect 464 112 465 113
rect 465 112 466 113
rect 466 112 467 113
rect 467 112 468 113
rect 468 112 469 113
rect 469 112 470 113
rect 470 112 471 113
rect 471 112 472 113
rect 472 112 473 113
rect 132 111 133 112
rect 133 111 134 112
rect 134 111 135 112
rect 135 111 136 112
rect 136 111 137 112
rect 137 111 138 112
rect 138 111 139 112
rect 139 111 140 112
rect 140 111 141 112
rect 141 111 142 112
rect 142 111 143 112
rect 143 111 144 112
rect 144 111 145 112
rect 145 111 146 112
rect 146 111 147 112
rect 147 111 148 112
rect 328 111 329 112
rect 329 111 330 112
rect 330 111 331 112
rect 331 111 332 112
rect 332 111 333 112
rect 333 111 334 112
rect 334 111 335 112
rect 335 111 336 112
rect 336 111 337 112
rect 337 111 338 112
rect 338 111 339 112
rect 339 111 340 112
rect 340 111 341 112
rect 341 111 342 112
rect 342 111 343 112
rect 343 111 344 112
rect 344 111 345 112
rect 345 111 346 112
rect 346 111 347 112
rect 347 111 348 112
rect 348 111 349 112
rect 349 111 350 112
rect 350 111 351 112
rect 351 111 352 112
rect 352 111 353 112
rect 353 111 354 112
rect 446 111 447 112
rect 447 111 448 112
rect 448 111 449 112
rect 449 111 450 112
rect 450 111 451 112
rect 451 111 452 112
rect 452 111 453 112
rect 453 111 454 112
rect 454 111 455 112
rect 455 111 456 112
rect 456 111 457 112
rect 457 111 458 112
rect 458 111 459 112
rect 459 111 460 112
rect 460 111 461 112
rect 461 111 462 112
rect 462 111 463 112
rect 463 111 464 112
rect 464 111 465 112
rect 465 111 466 112
rect 466 111 467 112
rect 467 111 468 112
rect 468 111 469 112
rect 469 111 470 112
rect 470 111 471 112
rect 471 111 472 112
rect 472 111 473 112
rect 132 110 133 111
rect 133 110 134 111
rect 134 110 135 111
rect 135 110 136 111
rect 136 110 137 111
rect 137 110 138 111
rect 138 110 139 111
rect 139 110 140 111
rect 140 110 141 111
rect 141 110 142 111
rect 142 110 143 111
rect 143 110 144 111
rect 144 110 145 111
rect 145 110 146 111
rect 146 110 147 111
rect 147 110 148 111
rect 328 110 329 111
rect 329 110 330 111
rect 330 110 331 111
rect 331 110 332 111
rect 332 110 333 111
rect 333 110 334 111
rect 334 110 335 111
rect 335 110 336 111
rect 336 110 337 111
rect 337 110 338 111
rect 338 110 339 111
rect 339 110 340 111
rect 340 110 341 111
rect 341 110 342 111
rect 342 110 343 111
rect 343 110 344 111
rect 344 110 345 111
rect 345 110 346 111
rect 346 110 347 111
rect 347 110 348 111
rect 348 110 349 111
rect 349 110 350 111
rect 350 110 351 111
rect 351 110 352 111
rect 352 110 353 111
rect 353 110 354 111
rect 446 110 447 111
rect 447 110 448 111
rect 448 110 449 111
rect 449 110 450 111
rect 450 110 451 111
rect 451 110 452 111
rect 452 110 453 111
rect 453 110 454 111
rect 454 110 455 111
rect 455 110 456 111
rect 456 110 457 111
rect 457 110 458 111
rect 458 110 459 111
rect 459 110 460 111
rect 460 110 461 111
rect 461 110 462 111
rect 462 110 463 111
rect 463 110 464 111
rect 464 110 465 111
rect 465 110 466 111
rect 466 110 467 111
rect 467 110 468 111
rect 468 110 469 111
rect 469 110 470 111
rect 470 110 471 111
rect 471 110 472 111
rect 132 109 133 110
rect 133 109 134 110
rect 134 109 135 110
rect 135 109 136 110
rect 136 109 137 110
rect 137 109 138 110
rect 138 109 139 110
rect 139 109 140 110
rect 140 109 141 110
rect 141 109 142 110
rect 142 109 143 110
rect 143 109 144 110
rect 144 109 145 110
rect 145 109 146 110
rect 146 109 147 110
rect 147 109 148 110
rect 148 109 149 110
rect 328 109 329 110
rect 329 109 330 110
rect 330 109 331 110
rect 331 109 332 110
rect 332 109 333 110
rect 333 109 334 110
rect 334 109 335 110
rect 335 109 336 110
rect 336 109 337 110
rect 337 109 338 110
rect 338 109 339 110
rect 339 109 340 110
rect 340 109 341 110
rect 341 109 342 110
rect 342 109 343 110
rect 343 109 344 110
rect 344 109 345 110
rect 345 109 346 110
rect 346 109 347 110
rect 347 109 348 110
rect 348 109 349 110
rect 349 109 350 110
rect 350 109 351 110
rect 351 109 352 110
rect 352 109 353 110
rect 353 109 354 110
rect 444 109 445 110
rect 445 109 446 110
rect 446 109 447 110
rect 447 109 448 110
rect 448 109 449 110
rect 449 109 450 110
rect 450 109 451 110
rect 451 109 452 110
rect 452 109 453 110
rect 453 109 454 110
rect 454 109 455 110
rect 455 109 456 110
rect 456 109 457 110
rect 457 109 458 110
rect 458 109 459 110
rect 459 109 460 110
rect 460 109 461 110
rect 461 109 462 110
rect 462 109 463 110
rect 463 109 464 110
rect 464 109 465 110
rect 465 109 466 110
rect 466 109 467 110
rect 467 109 468 110
rect 468 109 469 110
rect 469 109 470 110
rect 470 109 471 110
rect 471 109 472 110
rect 133 108 134 109
rect 134 108 135 109
rect 135 108 136 109
rect 136 108 137 109
rect 137 108 138 109
rect 138 108 139 109
rect 139 108 140 109
rect 140 108 141 109
rect 141 108 142 109
rect 142 108 143 109
rect 143 108 144 109
rect 144 108 145 109
rect 145 108 146 109
rect 146 108 147 109
rect 147 108 148 109
rect 148 108 149 109
rect 444 108 445 109
rect 445 108 446 109
rect 446 108 447 109
rect 447 108 448 109
rect 448 108 449 109
rect 449 108 450 109
rect 450 108 451 109
rect 451 108 452 109
rect 452 108 453 109
rect 453 108 454 109
rect 454 108 455 109
rect 455 108 456 109
rect 456 108 457 109
rect 457 108 458 109
rect 458 108 459 109
rect 459 108 460 109
rect 460 108 461 109
rect 461 108 462 109
rect 462 108 463 109
rect 463 108 464 109
rect 464 108 465 109
rect 465 108 466 109
rect 466 108 467 109
rect 467 108 468 109
rect 133 107 134 108
rect 134 107 135 108
rect 135 107 136 108
rect 136 107 137 108
rect 137 107 138 108
rect 138 107 139 108
rect 139 107 140 108
rect 140 107 141 108
rect 141 107 142 108
rect 142 107 143 108
rect 143 107 144 108
rect 144 107 145 108
rect 145 107 146 108
rect 146 107 147 108
rect 147 107 148 108
rect 148 107 149 108
rect 442 107 443 108
rect 443 107 444 108
rect 444 107 445 108
rect 445 107 446 108
rect 446 107 447 108
rect 447 107 448 108
rect 448 107 449 108
rect 449 107 450 108
rect 450 107 451 108
rect 451 107 452 108
rect 452 107 453 108
rect 453 107 454 108
rect 454 107 455 108
rect 455 107 456 108
rect 456 107 457 108
rect 457 107 458 108
rect 458 107 459 108
rect 459 107 460 108
rect 460 107 461 108
rect 461 107 462 108
rect 462 107 463 108
rect 463 107 464 108
rect 464 107 465 108
rect 465 107 466 108
rect 466 107 467 108
rect 467 107 468 108
rect 135 106 136 107
rect 136 106 137 107
rect 137 106 138 107
rect 138 106 139 107
rect 139 106 140 107
rect 140 106 141 107
rect 141 106 142 107
rect 142 106 143 107
rect 143 106 144 107
rect 144 106 145 107
rect 145 106 146 107
rect 146 106 147 107
rect 147 106 148 107
rect 148 106 149 107
rect 442 106 443 107
rect 443 106 444 107
rect 444 106 445 107
rect 445 106 446 107
rect 446 106 447 107
rect 447 106 448 107
rect 448 106 449 107
rect 449 106 450 107
rect 450 106 451 107
rect 451 106 452 107
rect 452 106 453 107
rect 453 106 454 107
rect 454 106 455 107
rect 455 106 456 107
rect 456 106 457 107
rect 457 106 458 107
rect 458 106 459 107
rect 459 106 460 107
rect 460 106 461 107
rect 461 106 462 107
rect 462 106 463 107
rect 463 106 464 107
rect 464 106 465 107
rect 465 106 466 107
rect 135 105 136 106
rect 136 105 137 106
rect 137 105 138 106
rect 138 105 139 106
rect 139 105 140 106
rect 140 105 141 106
rect 141 105 142 106
rect 142 105 143 106
rect 143 105 144 106
rect 144 105 145 106
rect 145 105 146 106
rect 146 105 147 106
rect 147 105 148 106
rect 148 105 149 106
rect 149 105 150 106
rect 150 105 151 106
rect 441 105 442 106
rect 442 105 443 106
rect 443 105 444 106
rect 444 105 445 106
rect 445 105 446 106
rect 446 105 447 106
rect 447 105 448 106
rect 448 105 449 106
rect 449 105 450 106
rect 450 105 451 106
rect 451 105 452 106
rect 452 105 453 106
rect 453 105 454 106
rect 454 105 455 106
rect 455 105 456 106
rect 456 105 457 106
rect 457 105 458 106
rect 458 105 459 106
rect 459 105 460 106
rect 460 105 461 106
rect 461 105 462 106
rect 462 105 463 106
rect 463 105 464 106
rect 464 105 465 106
rect 465 105 466 106
rect 137 104 138 105
rect 138 104 139 105
rect 139 104 140 105
rect 140 104 141 105
rect 141 104 142 105
rect 142 104 143 105
rect 143 104 144 105
rect 144 104 145 105
rect 145 104 146 105
rect 146 104 147 105
rect 147 104 148 105
rect 148 104 149 105
rect 149 104 150 105
rect 150 104 151 105
rect 441 104 442 105
rect 442 104 443 105
rect 443 104 444 105
rect 444 104 445 105
rect 445 104 446 105
rect 446 104 447 105
rect 447 104 448 105
rect 448 104 449 105
rect 449 104 450 105
rect 450 104 451 105
rect 451 104 452 105
rect 452 104 453 105
rect 453 104 454 105
rect 454 104 455 105
rect 455 104 456 105
rect 456 104 457 105
rect 457 104 458 105
rect 458 104 459 105
rect 459 104 460 105
rect 460 104 461 105
rect 461 104 462 105
rect 462 104 463 105
rect 463 104 464 105
rect 137 103 138 104
rect 138 103 139 104
rect 139 103 140 104
rect 140 103 141 104
rect 141 103 142 104
rect 142 103 143 104
rect 143 103 144 104
rect 144 103 145 104
rect 145 103 146 104
rect 146 103 147 104
rect 147 103 148 104
rect 148 103 149 104
rect 149 103 150 104
rect 150 103 151 104
rect 151 103 152 104
rect 152 103 153 104
rect 437 103 438 104
rect 438 103 439 104
rect 439 103 440 104
rect 440 103 441 104
rect 441 103 442 104
rect 442 103 443 104
rect 443 103 444 104
rect 444 103 445 104
rect 445 103 446 104
rect 446 103 447 104
rect 447 103 448 104
rect 448 103 449 104
rect 449 103 450 104
rect 450 103 451 104
rect 451 103 452 104
rect 452 103 453 104
rect 453 103 454 104
rect 454 103 455 104
rect 455 103 456 104
rect 456 103 457 104
rect 457 103 458 104
rect 458 103 459 104
rect 459 103 460 104
rect 460 103 461 104
rect 461 103 462 104
rect 462 103 463 104
rect 463 103 464 104
rect 139 102 140 103
rect 140 102 141 103
rect 141 102 142 103
rect 142 102 143 103
rect 143 102 144 103
rect 144 102 145 103
rect 145 102 146 103
rect 146 102 147 103
rect 147 102 148 103
rect 148 102 149 103
rect 149 102 150 103
rect 150 102 151 103
rect 151 102 152 103
rect 152 102 153 103
rect 437 102 438 103
rect 438 102 439 103
rect 439 102 440 103
rect 440 102 441 103
rect 441 102 442 103
rect 442 102 443 103
rect 443 102 444 103
rect 444 102 445 103
rect 445 102 446 103
rect 446 102 447 103
rect 447 102 448 103
rect 448 102 449 103
rect 449 102 450 103
rect 450 102 451 103
rect 451 102 452 103
rect 452 102 453 103
rect 453 102 454 103
rect 454 102 455 103
rect 455 102 456 103
rect 456 102 457 103
rect 457 102 458 103
rect 458 102 459 103
rect 459 102 460 103
rect 460 102 461 103
rect 461 102 462 103
rect 139 101 140 102
rect 140 101 141 102
rect 141 101 142 102
rect 142 101 143 102
rect 143 101 144 102
rect 144 101 145 102
rect 145 101 146 102
rect 146 101 147 102
rect 147 101 148 102
rect 148 101 149 102
rect 149 101 150 102
rect 150 101 151 102
rect 151 101 152 102
rect 152 101 153 102
rect 153 101 154 102
rect 154 101 155 102
rect 437 101 438 102
rect 438 101 439 102
rect 439 101 440 102
rect 440 101 441 102
rect 441 101 442 102
rect 442 101 443 102
rect 443 101 444 102
rect 444 101 445 102
rect 445 101 446 102
rect 446 101 447 102
rect 447 101 448 102
rect 448 101 449 102
rect 449 101 450 102
rect 450 101 451 102
rect 451 101 452 102
rect 452 101 453 102
rect 453 101 454 102
rect 454 101 455 102
rect 455 101 456 102
rect 456 101 457 102
rect 457 101 458 102
rect 458 101 459 102
rect 459 101 460 102
rect 460 101 461 102
rect 461 101 462 102
rect 139 100 140 101
rect 140 100 141 101
rect 141 100 142 101
rect 142 100 143 101
rect 143 100 144 101
rect 144 100 145 101
rect 145 100 146 101
rect 146 100 147 101
rect 147 100 148 101
rect 148 100 149 101
rect 149 100 150 101
rect 150 100 151 101
rect 151 100 152 101
rect 152 100 153 101
rect 153 100 154 101
rect 154 100 155 101
rect 437 100 438 101
rect 438 100 439 101
rect 439 100 440 101
rect 440 100 441 101
rect 441 100 442 101
rect 442 100 443 101
rect 443 100 444 101
rect 444 100 445 101
rect 445 100 446 101
rect 446 100 447 101
rect 447 100 448 101
rect 448 100 449 101
rect 449 100 450 101
rect 450 100 451 101
rect 451 100 452 101
rect 452 100 453 101
rect 453 100 454 101
rect 454 100 455 101
rect 455 100 456 101
rect 456 100 457 101
rect 457 100 458 101
rect 139 99 140 100
rect 140 99 141 100
rect 141 99 142 100
rect 142 99 143 100
rect 143 99 144 100
rect 144 99 145 100
rect 145 99 146 100
rect 146 99 147 100
rect 147 99 148 100
rect 148 99 149 100
rect 149 99 150 100
rect 150 99 151 100
rect 151 99 152 100
rect 152 99 153 100
rect 153 99 154 100
rect 154 99 155 100
rect 155 99 156 100
rect 156 99 157 100
rect 433 99 434 100
rect 434 99 435 100
rect 435 99 436 100
rect 436 99 437 100
rect 437 99 438 100
rect 438 99 439 100
rect 439 99 440 100
rect 440 99 441 100
rect 441 99 442 100
rect 442 99 443 100
rect 443 99 444 100
rect 444 99 445 100
rect 445 99 446 100
rect 446 99 447 100
rect 447 99 448 100
rect 448 99 449 100
rect 449 99 450 100
rect 450 99 451 100
rect 451 99 452 100
rect 452 99 453 100
rect 453 99 454 100
rect 454 99 455 100
rect 455 99 456 100
rect 456 99 457 100
rect 457 99 458 100
rect 141 98 142 99
rect 142 98 143 99
rect 143 98 144 99
rect 144 98 145 99
rect 145 98 146 99
rect 146 98 147 99
rect 147 98 148 99
rect 148 98 149 99
rect 149 98 150 99
rect 150 98 151 99
rect 151 98 152 99
rect 152 98 153 99
rect 153 98 154 99
rect 154 98 155 99
rect 155 98 156 99
rect 156 98 157 99
rect 433 98 434 99
rect 434 98 435 99
rect 435 98 436 99
rect 436 98 437 99
rect 437 98 438 99
rect 438 98 439 99
rect 439 98 440 99
rect 440 98 441 99
rect 441 98 442 99
rect 442 98 443 99
rect 443 98 444 99
rect 444 98 445 99
rect 445 98 446 99
rect 446 98 447 99
rect 447 98 448 99
rect 448 98 449 99
rect 449 98 450 99
rect 450 98 451 99
rect 451 98 452 99
rect 452 98 453 99
rect 453 98 454 99
rect 454 98 455 99
rect 455 98 456 99
rect 456 98 457 99
rect 141 97 142 98
rect 142 97 143 98
rect 143 97 144 98
rect 144 97 145 98
rect 145 97 146 98
rect 146 97 147 98
rect 147 97 148 98
rect 148 97 149 98
rect 149 97 150 98
rect 150 97 151 98
rect 151 97 152 98
rect 152 97 153 98
rect 153 97 154 98
rect 154 97 155 98
rect 155 97 156 98
rect 156 97 157 98
rect 157 97 158 98
rect 158 97 159 98
rect 431 97 432 98
rect 432 97 433 98
rect 433 97 434 98
rect 434 97 435 98
rect 435 97 436 98
rect 436 97 437 98
rect 437 97 438 98
rect 438 97 439 98
rect 439 97 440 98
rect 440 97 441 98
rect 441 97 442 98
rect 442 97 443 98
rect 443 97 444 98
rect 444 97 445 98
rect 445 97 446 98
rect 446 97 447 98
rect 447 97 448 98
rect 448 97 449 98
rect 449 97 450 98
rect 450 97 451 98
rect 451 97 452 98
rect 452 97 453 98
rect 453 97 454 98
rect 454 97 455 98
rect 455 97 456 98
rect 456 97 457 98
rect 143 96 144 97
rect 144 96 145 97
rect 145 96 146 97
rect 146 96 147 97
rect 147 96 148 97
rect 148 96 149 97
rect 149 96 150 97
rect 150 96 151 97
rect 151 96 152 97
rect 152 96 153 97
rect 153 96 154 97
rect 154 96 155 97
rect 155 96 156 97
rect 156 96 157 97
rect 157 96 158 97
rect 158 96 159 97
rect 431 96 432 97
rect 432 96 433 97
rect 433 96 434 97
rect 434 96 435 97
rect 435 96 436 97
rect 436 96 437 97
rect 437 96 438 97
rect 438 96 439 97
rect 439 96 440 97
rect 440 96 441 97
rect 441 96 442 97
rect 442 96 443 97
rect 443 96 444 97
rect 444 96 445 97
rect 445 96 446 97
rect 446 96 447 97
rect 447 96 448 97
rect 448 96 449 97
rect 449 96 450 97
rect 450 96 451 97
rect 451 96 452 97
rect 452 96 453 97
rect 453 96 454 97
rect 454 96 455 97
rect 143 95 144 96
rect 144 95 145 96
rect 145 95 146 96
rect 146 95 147 96
rect 147 95 148 96
rect 148 95 149 96
rect 149 95 150 96
rect 150 95 151 96
rect 151 95 152 96
rect 152 95 153 96
rect 153 95 154 96
rect 154 95 155 96
rect 155 95 156 96
rect 156 95 157 96
rect 157 95 158 96
rect 158 95 159 96
rect 159 95 160 96
rect 160 95 161 96
rect 161 95 162 96
rect 162 95 163 96
rect 429 95 430 96
rect 430 95 431 96
rect 431 95 432 96
rect 432 95 433 96
rect 433 95 434 96
rect 434 95 435 96
rect 435 95 436 96
rect 436 95 437 96
rect 437 95 438 96
rect 438 95 439 96
rect 439 95 440 96
rect 440 95 441 96
rect 441 95 442 96
rect 442 95 443 96
rect 443 95 444 96
rect 444 95 445 96
rect 445 95 446 96
rect 446 95 447 96
rect 447 95 448 96
rect 448 95 449 96
rect 449 95 450 96
rect 450 95 451 96
rect 451 95 452 96
rect 452 95 453 96
rect 453 95 454 96
rect 454 95 455 96
rect 145 94 146 95
rect 146 94 147 95
rect 147 94 148 95
rect 148 94 149 95
rect 149 94 150 95
rect 150 94 151 95
rect 151 94 152 95
rect 152 94 153 95
rect 153 94 154 95
rect 154 94 155 95
rect 155 94 156 95
rect 156 94 157 95
rect 157 94 158 95
rect 158 94 159 95
rect 159 94 160 95
rect 160 94 161 95
rect 161 94 162 95
rect 162 94 163 95
rect 429 94 430 95
rect 430 94 431 95
rect 431 94 432 95
rect 432 94 433 95
rect 433 94 434 95
rect 434 94 435 95
rect 435 94 436 95
rect 436 94 437 95
rect 437 94 438 95
rect 438 94 439 95
rect 439 94 440 95
rect 440 94 441 95
rect 441 94 442 95
rect 442 94 443 95
rect 443 94 444 95
rect 444 94 445 95
rect 445 94 446 95
rect 446 94 447 95
rect 447 94 448 95
rect 448 94 449 95
rect 449 94 450 95
rect 450 94 451 95
rect 145 93 146 94
rect 146 93 147 94
rect 147 93 148 94
rect 148 93 149 94
rect 149 93 150 94
rect 150 93 151 94
rect 151 93 152 94
rect 152 93 153 94
rect 153 93 154 94
rect 154 93 155 94
rect 155 93 156 94
rect 156 93 157 94
rect 157 93 158 94
rect 158 93 159 94
rect 159 93 160 94
rect 160 93 161 94
rect 161 93 162 94
rect 162 93 163 94
rect 427 93 428 94
rect 428 93 429 94
rect 429 93 430 94
rect 430 93 431 94
rect 431 93 432 94
rect 432 93 433 94
rect 433 93 434 94
rect 434 93 435 94
rect 435 93 436 94
rect 436 93 437 94
rect 437 93 438 94
rect 438 93 439 94
rect 439 93 440 94
rect 440 93 441 94
rect 441 93 442 94
rect 442 93 443 94
rect 443 93 444 94
rect 444 93 445 94
rect 445 93 446 94
rect 446 93 447 94
rect 447 93 448 94
rect 448 93 449 94
rect 449 93 450 94
rect 450 93 451 94
rect 147 92 148 93
rect 148 92 149 93
rect 149 92 150 93
rect 150 92 151 93
rect 151 92 152 93
rect 152 92 153 93
rect 153 92 154 93
rect 154 92 155 93
rect 155 92 156 93
rect 156 92 157 93
rect 157 92 158 93
rect 158 92 159 93
rect 159 92 160 93
rect 160 92 161 93
rect 161 92 162 93
rect 162 92 163 93
rect 427 92 428 93
rect 428 92 429 93
rect 429 92 430 93
rect 430 92 431 93
rect 431 92 432 93
rect 432 92 433 93
rect 433 92 434 93
rect 434 92 435 93
rect 435 92 436 93
rect 436 92 437 93
rect 437 92 438 93
rect 438 92 439 93
rect 439 92 440 93
rect 440 92 441 93
rect 441 92 442 93
rect 442 92 443 93
rect 443 92 444 93
rect 444 92 445 93
rect 445 92 446 93
rect 446 92 447 93
rect 447 92 448 93
rect 448 92 449 93
rect 147 91 148 92
rect 148 91 149 92
rect 149 91 150 92
rect 150 91 151 92
rect 151 91 152 92
rect 152 91 153 92
rect 153 91 154 92
rect 154 91 155 92
rect 155 91 156 92
rect 156 91 157 92
rect 157 91 158 92
rect 158 91 159 92
rect 159 91 160 92
rect 160 91 161 92
rect 161 91 162 92
rect 162 91 163 92
rect 163 91 164 92
rect 164 91 165 92
rect 165 91 166 92
rect 426 91 427 92
rect 427 91 428 92
rect 428 91 429 92
rect 429 91 430 92
rect 430 91 431 92
rect 431 91 432 92
rect 432 91 433 92
rect 433 91 434 92
rect 434 91 435 92
rect 435 91 436 92
rect 436 91 437 92
rect 437 91 438 92
rect 438 91 439 92
rect 439 91 440 92
rect 440 91 441 92
rect 441 91 442 92
rect 442 91 443 92
rect 443 91 444 92
rect 444 91 445 92
rect 445 91 446 92
rect 446 91 447 92
rect 447 91 448 92
rect 448 91 449 92
rect 148 90 149 91
rect 149 90 150 91
rect 150 90 151 91
rect 151 90 152 91
rect 152 90 153 91
rect 153 90 154 91
rect 154 90 155 91
rect 155 90 156 91
rect 156 90 157 91
rect 157 90 158 91
rect 158 90 159 91
rect 159 90 160 91
rect 160 90 161 91
rect 161 90 162 91
rect 162 90 163 91
rect 163 90 164 91
rect 164 90 165 91
rect 165 90 166 91
rect 426 90 427 91
rect 427 90 428 91
rect 428 90 429 91
rect 429 90 430 91
rect 430 90 431 91
rect 431 90 432 91
rect 432 90 433 91
rect 433 90 434 91
rect 434 90 435 91
rect 435 90 436 91
rect 436 90 437 91
rect 437 90 438 91
rect 438 90 439 91
rect 439 90 440 91
rect 440 90 441 91
rect 441 90 442 91
rect 442 90 443 91
rect 443 90 444 91
rect 444 90 445 91
rect 445 90 446 91
rect 446 90 447 91
rect 148 89 149 90
rect 149 89 150 90
rect 150 89 151 90
rect 151 89 152 90
rect 152 89 153 90
rect 153 89 154 90
rect 154 89 155 90
rect 155 89 156 90
rect 156 89 157 90
rect 157 89 158 90
rect 158 89 159 90
rect 159 89 160 90
rect 160 89 161 90
rect 161 89 162 90
rect 162 89 163 90
rect 163 89 164 90
rect 164 89 165 90
rect 165 89 166 90
rect 166 89 167 90
rect 167 89 168 90
rect 424 89 425 90
rect 425 89 426 90
rect 426 89 427 90
rect 427 89 428 90
rect 428 89 429 90
rect 429 89 430 90
rect 430 89 431 90
rect 431 89 432 90
rect 432 89 433 90
rect 433 89 434 90
rect 434 89 435 90
rect 435 89 436 90
rect 436 89 437 90
rect 437 89 438 90
rect 438 89 439 90
rect 439 89 440 90
rect 440 89 441 90
rect 441 89 442 90
rect 442 89 443 90
rect 443 89 444 90
rect 444 89 445 90
rect 445 89 446 90
rect 446 89 447 90
rect 150 88 151 89
rect 151 88 152 89
rect 152 88 153 89
rect 153 88 154 89
rect 154 88 155 89
rect 155 88 156 89
rect 156 88 157 89
rect 157 88 158 89
rect 158 88 159 89
rect 159 88 160 89
rect 160 88 161 89
rect 161 88 162 89
rect 162 88 163 89
rect 163 88 164 89
rect 164 88 165 89
rect 165 88 166 89
rect 166 88 167 89
rect 167 88 168 89
rect 424 88 425 89
rect 425 88 426 89
rect 426 88 427 89
rect 427 88 428 89
rect 428 88 429 89
rect 429 88 430 89
rect 430 88 431 89
rect 431 88 432 89
rect 432 88 433 89
rect 433 88 434 89
rect 434 88 435 89
rect 435 88 436 89
rect 436 88 437 89
rect 437 88 438 89
rect 438 88 439 89
rect 439 88 440 89
rect 440 88 441 89
rect 441 88 442 89
rect 442 88 443 89
rect 150 87 151 88
rect 151 87 152 88
rect 152 87 153 88
rect 153 87 154 88
rect 154 87 155 88
rect 155 87 156 88
rect 156 87 157 88
rect 157 87 158 88
rect 158 87 159 88
rect 159 87 160 88
rect 160 87 161 88
rect 161 87 162 88
rect 162 87 163 88
rect 163 87 164 88
rect 164 87 165 88
rect 165 87 166 88
rect 166 87 167 88
rect 167 87 168 88
rect 168 87 169 88
rect 169 87 170 88
rect 422 87 423 88
rect 423 87 424 88
rect 424 87 425 88
rect 425 87 426 88
rect 426 87 427 88
rect 427 87 428 88
rect 428 87 429 88
rect 429 87 430 88
rect 430 87 431 88
rect 431 87 432 88
rect 432 87 433 88
rect 433 87 434 88
rect 434 87 435 88
rect 435 87 436 88
rect 436 87 437 88
rect 437 87 438 88
rect 438 87 439 88
rect 439 87 440 88
rect 440 87 441 88
rect 441 87 442 88
rect 442 87 443 88
rect 152 86 153 87
rect 153 86 154 87
rect 154 86 155 87
rect 155 86 156 87
rect 156 86 157 87
rect 157 86 158 87
rect 158 86 159 87
rect 159 86 160 87
rect 160 86 161 87
rect 161 86 162 87
rect 162 86 163 87
rect 163 86 164 87
rect 164 86 165 87
rect 165 86 166 87
rect 166 86 167 87
rect 167 86 168 87
rect 168 86 169 87
rect 169 86 170 87
rect 422 86 423 87
rect 423 86 424 87
rect 424 86 425 87
rect 425 86 426 87
rect 426 86 427 87
rect 427 86 428 87
rect 428 86 429 87
rect 429 86 430 87
rect 430 86 431 87
rect 431 86 432 87
rect 432 86 433 87
rect 433 86 434 87
rect 434 86 435 87
rect 435 86 436 87
rect 436 86 437 87
rect 437 86 438 87
rect 438 86 439 87
rect 439 86 440 87
rect 440 86 441 87
rect 441 86 442 87
rect 152 85 153 86
rect 153 85 154 86
rect 154 85 155 86
rect 155 85 156 86
rect 156 85 157 86
rect 157 85 158 86
rect 158 85 159 86
rect 159 85 160 86
rect 160 85 161 86
rect 161 85 162 86
rect 162 85 163 86
rect 163 85 164 86
rect 164 85 165 86
rect 165 85 166 86
rect 166 85 167 86
rect 167 85 168 86
rect 168 85 169 86
rect 169 85 170 86
rect 170 85 171 86
rect 171 85 172 86
rect 420 85 421 86
rect 421 85 422 86
rect 422 85 423 86
rect 423 85 424 86
rect 424 85 425 86
rect 425 85 426 86
rect 426 85 427 86
rect 427 85 428 86
rect 428 85 429 86
rect 429 85 430 86
rect 430 85 431 86
rect 431 85 432 86
rect 432 85 433 86
rect 433 85 434 86
rect 434 85 435 86
rect 435 85 436 86
rect 436 85 437 86
rect 437 85 438 86
rect 438 85 439 86
rect 439 85 440 86
rect 440 85 441 86
rect 441 85 442 86
rect 154 84 155 85
rect 155 84 156 85
rect 156 84 157 85
rect 157 84 158 85
rect 158 84 159 85
rect 159 84 160 85
rect 160 84 161 85
rect 161 84 162 85
rect 162 84 163 85
rect 163 84 164 85
rect 164 84 165 85
rect 165 84 166 85
rect 166 84 167 85
rect 167 84 168 85
rect 168 84 169 85
rect 169 84 170 85
rect 170 84 171 85
rect 171 84 172 85
rect 420 84 421 85
rect 421 84 422 85
rect 422 84 423 85
rect 423 84 424 85
rect 424 84 425 85
rect 425 84 426 85
rect 426 84 427 85
rect 427 84 428 85
rect 428 84 429 85
rect 429 84 430 85
rect 430 84 431 85
rect 431 84 432 85
rect 432 84 433 85
rect 433 84 434 85
rect 434 84 435 85
rect 435 84 436 85
rect 436 84 437 85
rect 437 84 438 85
rect 438 84 439 85
rect 439 84 440 85
rect 154 83 155 84
rect 155 83 156 84
rect 156 83 157 84
rect 157 83 158 84
rect 158 83 159 84
rect 159 83 160 84
rect 160 83 161 84
rect 161 83 162 84
rect 162 83 163 84
rect 163 83 164 84
rect 164 83 165 84
rect 165 83 166 84
rect 166 83 167 84
rect 167 83 168 84
rect 168 83 169 84
rect 169 83 170 84
rect 170 83 171 84
rect 171 83 172 84
rect 172 83 173 84
rect 173 83 174 84
rect 418 83 419 84
rect 419 83 420 84
rect 420 83 421 84
rect 421 83 422 84
rect 422 83 423 84
rect 423 83 424 84
rect 424 83 425 84
rect 425 83 426 84
rect 426 83 427 84
rect 427 83 428 84
rect 428 83 429 84
rect 429 83 430 84
rect 430 83 431 84
rect 431 83 432 84
rect 432 83 433 84
rect 433 83 434 84
rect 434 83 435 84
rect 435 83 436 84
rect 436 83 437 84
rect 437 83 438 84
rect 438 83 439 84
rect 439 83 440 84
rect 156 82 157 83
rect 157 82 158 83
rect 158 82 159 83
rect 159 82 160 83
rect 160 82 161 83
rect 161 82 162 83
rect 162 82 163 83
rect 163 82 164 83
rect 164 82 165 83
rect 165 82 166 83
rect 166 82 167 83
rect 167 82 168 83
rect 168 82 169 83
rect 169 82 170 83
rect 170 82 171 83
rect 171 82 172 83
rect 172 82 173 83
rect 173 82 174 83
rect 418 82 419 83
rect 419 82 420 83
rect 420 82 421 83
rect 421 82 422 83
rect 422 82 423 83
rect 423 82 424 83
rect 424 82 425 83
rect 425 82 426 83
rect 426 82 427 83
rect 427 82 428 83
rect 428 82 429 83
rect 429 82 430 83
rect 430 82 431 83
rect 431 82 432 83
rect 432 82 433 83
rect 433 82 434 83
rect 434 82 435 83
rect 435 82 436 83
rect 156 81 157 82
rect 157 81 158 82
rect 158 81 159 82
rect 159 81 160 82
rect 160 81 161 82
rect 161 81 162 82
rect 162 81 163 82
rect 163 81 164 82
rect 164 81 165 82
rect 165 81 166 82
rect 166 81 167 82
rect 167 81 168 82
rect 168 81 169 82
rect 169 81 170 82
rect 170 81 171 82
rect 171 81 172 82
rect 172 81 173 82
rect 173 81 174 82
rect 174 81 175 82
rect 175 81 176 82
rect 416 81 417 82
rect 417 81 418 82
rect 418 81 419 82
rect 419 81 420 82
rect 420 81 421 82
rect 421 81 422 82
rect 422 81 423 82
rect 423 81 424 82
rect 424 81 425 82
rect 425 81 426 82
rect 426 81 427 82
rect 427 81 428 82
rect 428 81 429 82
rect 429 81 430 82
rect 430 81 431 82
rect 431 81 432 82
rect 432 81 433 82
rect 433 81 434 82
rect 434 81 435 82
rect 435 81 436 82
rect 158 80 159 81
rect 159 80 160 81
rect 160 80 161 81
rect 161 80 162 81
rect 162 80 163 81
rect 163 80 164 81
rect 164 80 165 81
rect 165 80 166 81
rect 166 80 167 81
rect 167 80 168 81
rect 168 80 169 81
rect 169 80 170 81
rect 170 80 171 81
rect 171 80 172 81
rect 172 80 173 81
rect 173 80 174 81
rect 174 80 175 81
rect 175 80 176 81
rect 416 80 417 81
rect 417 80 418 81
rect 418 80 419 81
rect 419 80 420 81
rect 420 80 421 81
rect 421 80 422 81
rect 422 80 423 81
rect 423 80 424 81
rect 424 80 425 81
rect 425 80 426 81
rect 426 80 427 81
rect 427 80 428 81
rect 428 80 429 81
rect 429 80 430 81
rect 430 80 431 81
rect 431 80 432 81
rect 432 80 433 81
rect 433 80 434 81
rect 158 79 159 80
rect 159 79 160 80
rect 160 79 161 80
rect 161 79 162 80
rect 162 79 163 80
rect 163 79 164 80
rect 164 79 165 80
rect 165 79 166 80
rect 166 79 167 80
rect 167 79 168 80
rect 168 79 169 80
rect 169 79 170 80
rect 170 79 171 80
rect 171 79 172 80
rect 172 79 173 80
rect 173 79 174 80
rect 174 79 175 80
rect 175 79 176 80
rect 176 79 177 80
rect 177 79 178 80
rect 178 79 179 80
rect 414 79 415 80
rect 415 79 416 80
rect 416 79 417 80
rect 417 79 418 80
rect 418 79 419 80
rect 419 79 420 80
rect 420 79 421 80
rect 421 79 422 80
rect 422 79 423 80
rect 423 79 424 80
rect 424 79 425 80
rect 425 79 426 80
rect 426 79 427 80
rect 427 79 428 80
rect 428 79 429 80
rect 429 79 430 80
rect 430 79 431 80
rect 431 79 432 80
rect 432 79 433 80
rect 433 79 434 80
rect 162 78 163 79
rect 163 78 164 79
rect 164 78 165 79
rect 165 78 166 79
rect 166 78 167 79
rect 167 78 168 79
rect 168 78 169 79
rect 169 78 170 79
rect 170 78 171 79
rect 171 78 172 79
rect 172 78 173 79
rect 173 78 174 79
rect 174 78 175 79
rect 175 78 176 79
rect 176 78 177 79
rect 177 78 178 79
rect 178 78 179 79
rect 414 78 415 79
rect 415 78 416 79
rect 416 78 417 79
rect 417 78 418 79
rect 418 78 419 79
rect 419 78 420 79
rect 420 78 421 79
rect 421 78 422 79
rect 422 78 423 79
rect 423 78 424 79
rect 424 78 425 79
rect 425 78 426 79
rect 426 78 427 79
rect 427 78 428 79
rect 428 78 429 79
rect 429 78 430 79
rect 162 77 163 78
rect 163 77 164 78
rect 164 77 165 78
rect 165 77 166 78
rect 166 77 167 78
rect 167 77 168 78
rect 168 77 169 78
rect 169 77 170 78
rect 170 77 171 78
rect 171 77 172 78
rect 172 77 173 78
rect 173 77 174 78
rect 174 77 175 78
rect 175 77 176 78
rect 176 77 177 78
rect 177 77 178 78
rect 178 77 179 78
rect 414 77 415 78
rect 415 77 416 78
rect 416 77 417 78
rect 417 77 418 78
rect 418 77 419 78
rect 419 77 420 78
rect 420 77 421 78
rect 421 77 422 78
rect 422 77 423 78
rect 423 77 424 78
rect 424 77 425 78
rect 425 77 426 78
rect 426 77 427 78
rect 427 77 428 78
rect 428 77 429 78
rect 429 77 430 78
rect 162 76 163 77
rect 163 76 164 77
rect 164 76 165 77
rect 165 76 166 77
rect 166 76 167 77
rect 167 76 168 77
rect 168 76 169 77
rect 169 76 170 77
rect 170 76 171 77
rect 171 76 172 77
rect 172 76 173 77
rect 173 76 174 77
rect 174 76 175 77
rect 175 76 176 77
rect 176 76 177 77
rect 177 76 178 77
rect 178 76 179 77
rect 179 76 180 77
rect 180 76 181 77
rect 411 76 412 77
rect 412 76 413 77
rect 413 76 414 77
rect 414 76 415 77
rect 415 76 416 77
rect 416 76 417 77
rect 417 76 418 77
rect 418 76 419 77
rect 419 76 420 77
rect 420 76 421 77
rect 421 76 422 77
rect 422 76 423 77
rect 423 76 424 77
rect 424 76 425 77
rect 425 76 426 77
rect 426 76 427 77
rect 427 76 428 77
rect 428 76 429 77
rect 429 76 430 77
rect 162 75 163 76
rect 163 75 164 76
rect 164 75 165 76
rect 165 75 166 76
rect 166 75 167 76
rect 167 75 168 76
rect 168 75 169 76
rect 169 75 170 76
rect 170 75 171 76
rect 171 75 172 76
rect 172 75 173 76
rect 173 75 174 76
rect 174 75 175 76
rect 175 75 176 76
rect 176 75 177 76
rect 177 75 178 76
rect 178 75 179 76
rect 179 75 180 76
rect 180 75 181 76
rect 411 75 412 76
rect 412 75 413 76
rect 413 75 414 76
rect 414 75 415 76
rect 415 75 416 76
rect 416 75 417 76
rect 417 75 418 76
rect 418 75 419 76
rect 419 75 420 76
rect 420 75 421 76
rect 421 75 422 76
rect 422 75 423 76
rect 423 75 424 76
rect 424 75 425 76
rect 425 75 426 76
rect 426 75 427 76
rect 427 75 428 76
rect 162 74 163 75
rect 163 74 164 75
rect 164 74 165 75
rect 165 74 166 75
rect 166 74 167 75
rect 167 74 168 75
rect 168 74 169 75
rect 169 74 170 75
rect 170 74 171 75
rect 171 74 172 75
rect 172 74 173 75
rect 173 74 174 75
rect 174 74 175 75
rect 175 74 176 75
rect 176 74 177 75
rect 177 74 178 75
rect 178 74 179 75
rect 179 74 180 75
rect 180 74 181 75
rect 181 74 182 75
rect 182 74 183 75
rect 183 74 184 75
rect 184 74 185 75
rect 409 74 410 75
rect 410 74 411 75
rect 411 74 412 75
rect 412 74 413 75
rect 413 74 414 75
rect 414 74 415 75
rect 415 74 416 75
rect 416 74 417 75
rect 417 74 418 75
rect 418 74 419 75
rect 419 74 420 75
rect 420 74 421 75
rect 421 74 422 75
rect 422 74 423 75
rect 423 74 424 75
rect 424 74 425 75
rect 425 74 426 75
rect 426 74 427 75
rect 427 74 428 75
rect 165 73 166 74
rect 166 73 167 74
rect 167 73 168 74
rect 168 73 169 74
rect 169 73 170 74
rect 170 73 171 74
rect 171 73 172 74
rect 172 73 173 74
rect 173 73 174 74
rect 174 73 175 74
rect 175 73 176 74
rect 176 73 177 74
rect 177 73 178 74
rect 178 73 179 74
rect 179 73 180 74
rect 180 73 181 74
rect 181 73 182 74
rect 182 73 183 74
rect 183 73 184 74
rect 184 73 185 74
rect 409 73 410 74
rect 410 73 411 74
rect 411 73 412 74
rect 412 73 413 74
rect 413 73 414 74
rect 414 73 415 74
rect 415 73 416 74
rect 416 73 417 74
rect 417 73 418 74
rect 418 73 419 74
rect 419 73 420 74
rect 420 73 421 74
rect 421 73 422 74
rect 422 73 423 74
rect 423 73 424 74
rect 424 73 425 74
rect 165 72 166 73
rect 166 72 167 73
rect 167 72 168 73
rect 168 72 169 73
rect 169 72 170 73
rect 170 72 171 73
rect 171 72 172 73
rect 172 72 173 73
rect 173 72 174 73
rect 174 72 175 73
rect 175 72 176 73
rect 176 72 177 73
rect 177 72 178 73
rect 178 72 179 73
rect 179 72 180 73
rect 180 72 181 73
rect 181 72 182 73
rect 182 72 183 73
rect 183 72 184 73
rect 184 72 185 73
rect 185 72 186 73
rect 186 72 187 73
rect 407 72 408 73
rect 408 72 409 73
rect 409 72 410 73
rect 410 72 411 73
rect 411 72 412 73
rect 412 72 413 73
rect 413 72 414 73
rect 414 72 415 73
rect 415 72 416 73
rect 416 72 417 73
rect 417 72 418 73
rect 418 72 419 73
rect 419 72 420 73
rect 420 72 421 73
rect 421 72 422 73
rect 422 72 423 73
rect 423 72 424 73
rect 424 72 425 73
rect 167 71 168 72
rect 168 71 169 72
rect 169 71 170 72
rect 170 71 171 72
rect 171 71 172 72
rect 172 71 173 72
rect 173 71 174 72
rect 174 71 175 72
rect 175 71 176 72
rect 176 71 177 72
rect 177 71 178 72
rect 178 71 179 72
rect 179 71 180 72
rect 180 71 181 72
rect 181 71 182 72
rect 182 71 183 72
rect 183 71 184 72
rect 184 71 185 72
rect 185 71 186 72
rect 186 71 187 72
rect 407 71 408 72
rect 408 71 409 72
rect 409 71 410 72
rect 410 71 411 72
rect 411 71 412 72
rect 412 71 413 72
rect 413 71 414 72
rect 414 71 415 72
rect 415 71 416 72
rect 416 71 417 72
rect 417 71 418 72
rect 418 71 419 72
rect 419 71 420 72
rect 420 71 421 72
rect 421 71 422 72
rect 422 71 423 72
rect 167 70 168 71
rect 168 70 169 71
rect 169 70 170 71
rect 170 70 171 71
rect 171 70 172 71
rect 172 70 173 71
rect 173 70 174 71
rect 174 70 175 71
rect 175 70 176 71
rect 176 70 177 71
rect 177 70 178 71
rect 178 70 179 71
rect 179 70 180 71
rect 180 70 181 71
rect 181 70 182 71
rect 182 70 183 71
rect 183 70 184 71
rect 184 70 185 71
rect 185 70 186 71
rect 186 70 187 71
rect 187 70 188 71
rect 188 70 189 71
rect 405 70 406 71
rect 406 70 407 71
rect 407 70 408 71
rect 408 70 409 71
rect 409 70 410 71
rect 410 70 411 71
rect 411 70 412 71
rect 412 70 413 71
rect 413 70 414 71
rect 414 70 415 71
rect 415 70 416 71
rect 416 70 417 71
rect 417 70 418 71
rect 418 70 419 71
rect 419 70 420 71
rect 420 70 421 71
rect 421 70 422 71
rect 422 70 423 71
rect 169 69 170 70
rect 170 69 171 70
rect 171 69 172 70
rect 172 69 173 70
rect 173 69 174 70
rect 174 69 175 70
rect 175 69 176 70
rect 176 69 177 70
rect 177 69 178 70
rect 178 69 179 70
rect 179 69 180 70
rect 180 69 181 70
rect 181 69 182 70
rect 182 69 183 70
rect 183 69 184 70
rect 184 69 185 70
rect 185 69 186 70
rect 186 69 187 70
rect 187 69 188 70
rect 188 69 189 70
rect 405 69 406 70
rect 406 69 407 70
rect 407 69 408 70
rect 408 69 409 70
rect 409 69 410 70
rect 410 69 411 70
rect 411 69 412 70
rect 412 69 413 70
rect 413 69 414 70
rect 414 69 415 70
rect 415 69 416 70
rect 416 69 417 70
rect 417 69 418 70
rect 418 69 419 70
rect 169 68 170 69
rect 170 68 171 69
rect 171 68 172 69
rect 172 68 173 69
rect 173 68 174 69
rect 174 68 175 69
rect 175 68 176 69
rect 176 68 177 69
rect 177 68 178 69
rect 178 68 179 69
rect 179 68 180 69
rect 180 68 181 69
rect 181 68 182 69
rect 182 68 183 69
rect 183 68 184 69
rect 184 68 185 69
rect 185 68 186 69
rect 186 68 187 69
rect 187 68 188 69
rect 188 68 189 69
rect 189 68 190 69
rect 190 68 191 69
rect 191 68 192 69
rect 403 68 404 69
rect 404 68 405 69
rect 405 68 406 69
rect 406 68 407 69
rect 407 68 408 69
rect 408 68 409 69
rect 409 68 410 69
rect 410 68 411 69
rect 411 68 412 69
rect 412 68 413 69
rect 413 68 414 69
rect 414 68 415 69
rect 415 68 416 69
rect 416 68 417 69
rect 417 68 418 69
rect 418 68 419 69
rect 171 67 172 68
rect 172 67 173 68
rect 173 67 174 68
rect 174 67 175 68
rect 175 67 176 68
rect 176 67 177 68
rect 177 67 178 68
rect 178 67 179 68
rect 179 67 180 68
rect 180 67 181 68
rect 181 67 182 68
rect 182 67 183 68
rect 183 67 184 68
rect 184 67 185 68
rect 185 67 186 68
rect 186 67 187 68
rect 187 67 188 68
rect 188 67 189 68
rect 189 67 190 68
rect 190 67 191 68
rect 191 67 192 68
rect 403 67 404 68
rect 404 67 405 68
rect 405 67 406 68
rect 406 67 407 68
rect 407 67 408 68
rect 408 67 409 68
rect 409 67 410 68
rect 410 67 411 68
rect 411 67 412 68
rect 412 67 413 68
rect 413 67 414 68
rect 414 67 415 68
rect 415 67 416 68
rect 416 67 417 68
rect 171 66 172 67
rect 172 66 173 67
rect 173 66 174 67
rect 174 66 175 67
rect 175 66 176 67
rect 176 66 177 67
rect 177 66 178 67
rect 178 66 179 67
rect 179 66 180 67
rect 180 66 181 67
rect 181 66 182 67
rect 182 66 183 67
rect 183 66 184 67
rect 184 66 185 67
rect 185 66 186 67
rect 186 66 187 67
rect 187 66 188 67
rect 188 66 189 67
rect 189 66 190 67
rect 190 66 191 67
rect 191 66 192 67
rect 192 66 193 67
rect 193 66 194 67
rect 194 66 195 67
rect 195 66 196 67
rect 401 66 402 67
rect 402 66 403 67
rect 403 66 404 67
rect 404 66 405 67
rect 405 66 406 67
rect 406 66 407 67
rect 407 66 408 67
rect 408 66 409 67
rect 409 66 410 67
rect 410 66 411 67
rect 411 66 412 67
rect 412 66 413 67
rect 413 66 414 67
rect 414 66 415 67
rect 415 66 416 67
rect 416 66 417 67
rect 175 65 176 66
rect 176 65 177 66
rect 177 65 178 66
rect 178 65 179 66
rect 179 65 180 66
rect 180 65 181 66
rect 181 65 182 66
rect 182 65 183 66
rect 183 65 184 66
rect 184 65 185 66
rect 185 65 186 66
rect 186 65 187 66
rect 187 65 188 66
rect 188 65 189 66
rect 189 65 190 66
rect 190 65 191 66
rect 191 65 192 66
rect 192 65 193 66
rect 193 65 194 66
rect 194 65 195 66
rect 195 65 196 66
rect 401 65 402 66
rect 402 65 403 66
rect 403 65 404 66
rect 404 65 405 66
rect 405 65 406 66
rect 406 65 407 66
rect 407 65 408 66
rect 408 65 409 66
rect 409 65 410 66
rect 410 65 411 66
rect 411 65 412 66
rect 412 65 413 66
rect 175 64 176 65
rect 176 64 177 65
rect 177 64 178 65
rect 178 64 179 65
rect 179 64 180 65
rect 180 64 181 65
rect 181 64 182 65
rect 182 64 183 65
rect 183 64 184 65
rect 184 64 185 65
rect 185 64 186 65
rect 186 64 187 65
rect 187 64 188 65
rect 188 64 189 65
rect 189 64 190 65
rect 190 64 191 65
rect 191 64 192 65
rect 192 64 193 65
rect 193 64 194 65
rect 194 64 195 65
rect 195 64 196 65
rect 196 64 197 65
rect 197 64 198 65
rect 397 64 398 65
rect 398 64 399 65
rect 399 64 400 65
rect 400 64 401 65
rect 401 64 402 65
rect 402 64 403 65
rect 403 64 404 65
rect 404 64 405 65
rect 405 64 406 65
rect 406 64 407 65
rect 407 64 408 65
rect 408 64 409 65
rect 409 64 410 65
rect 410 64 411 65
rect 411 64 412 65
rect 412 64 413 65
rect 176 63 177 64
rect 177 63 178 64
rect 178 63 179 64
rect 179 63 180 64
rect 180 63 181 64
rect 181 63 182 64
rect 182 63 183 64
rect 183 63 184 64
rect 184 63 185 64
rect 185 63 186 64
rect 186 63 187 64
rect 187 63 188 64
rect 188 63 189 64
rect 189 63 190 64
rect 190 63 191 64
rect 191 63 192 64
rect 192 63 193 64
rect 193 63 194 64
rect 194 63 195 64
rect 195 63 196 64
rect 196 63 197 64
rect 197 63 198 64
rect 397 63 398 64
rect 398 63 399 64
rect 399 63 400 64
rect 400 63 401 64
rect 401 63 402 64
rect 402 63 403 64
rect 403 63 404 64
rect 404 63 405 64
rect 405 63 406 64
rect 406 63 407 64
rect 407 63 408 64
rect 408 63 409 64
rect 409 63 410 64
rect 410 63 411 64
rect 411 63 412 64
rect 176 62 177 63
rect 177 62 178 63
rect 178 62 179 63
rect 179 62 180 63
rect 180 62 181 63
rect 181 62 182 63
rect 182 62 183 63
rect 183 62 184 63
rect 184 62 185 63
rect 185 62 186 63
rect 186 62 187 63
rect 187 62 188 63
rect 188 62 189 63
rect 189 62 190 63
rect 190 62 191 63
rect 191 62 192 63
rect 192 62 193 63
rect 193 62 194 63
rect 194 62 195 63
rect 195 62 196 63
rect 196 62 197 63
rect 197 62 198 63
rect 198 62 199 63
rect 199 62 200 63
rect 200 62 201 63
rect 201 62 202 63
rect 396 62 397 63
rect 397 62 398 63
rect 398 62 399 63
rect 399 62 400 63
rect 400 62 401 63
rect 401 62 402 63
rect 402 62 403 63
rect 403 62 404 63
rect 404 62 405 63
rect 405 62 406 63
rect 406 62 407 63
rect 407 62 408 63
rect 408 62 409 63
rect 409 62 410 63
rect 410 62 411 63
rect 411 62 412 63
rect 180 61 181 62
rect 181 61 182 62
rect 182 61 183 62
rect 183 61 184 62
rect 184 61 185 62
rect 185 61 186 62
rect 186 61 187 62
rect 187 61 188 62
rect 188 61 189 62
rect 189 61 190 62
rect 190 61 191 62
rect 191 61 192 62
rect 192 61 193 62
rect 193 61 194 62
rect 194 61 195 62
rect 195 61 196 62
rect 196 61 197 62
rect 197 61 198 62
rect 198 61 199 62
rect 199 61 200 62
rect 200 61 201 62
rect 201 61 202 62
rect 396 61 397 62
rect 397 61 398 62
rect 398 61 399 62
rect 399 61 400 62
rect 400 61 401 62
rect 401 61 402 62
rect 402 61 403 62
rect 403 61 404 62
rect 404 61 405 62
rect 405 61 406 62
rect 406 61 407 62
rect 407 61 408 62
rect 180 60 181 61
rect 181 60 182 61
rect 182 60 183 61
rect 183 60 184 61
rect 184 60 185 61
rect 185 60 186 61
rect 186 60 187 61
rect 187 60 188 61
rect 188 60 189 61
rect 189 60 190 61
rect 190 60 191 61
rect 191 60 192 61
rect 192 60 193 61
rect 193 60 194 61
rect 194 60 195 61
rect 195 60 196 61
rect 196 60 197 61
rect 197 60 198 61
rect 198 60 199 61
rect 199 60 200 61
rect 200 60 201 61
rect 201 60 202 61
rect 202 60 203 61
rect 203 60 204 61
rect 204 60 205 61
rect 205 60 206 61
rect 317 60 318 61
rect 318 60 319 61
rect 319 60 320 61
rect 320 60 321 61
rect 321 60 322 61
rect 322 60 323 61
rect 323 60 324 61
rect 394 60 395 61
rect 395 60 396 61
rect 396 60 397 61
rect 397 60 398 61
rect 398 60 399 61
rect 399 60 400 61
rect 400 60 401 61
rect 401 60 402 61
rect 402 60 403 61
rect 403 60 404 61
rect 404 60 405 61
rect 405 60 406 61
rect 406 60 407 61
rect 407 60 408 61
rect 182 59 183 60
rect 183 59 184 60
rect 184 59 185 60
rect 185 59 186 60
rect 186 59 187 60
rect 187 59 188 60
rect 188 59 189 60
rect 189 59 190 60
rect 190 59 191 60
rect 191 59 192 60
rect 192 59 193 60
rect 193 59 194 60
rect 194 59 195 60
rect 195 59 196 60
rect 196 59 197 60
rect 197 59 198 60
rect 198 59 199 60
rect 199 59 200 60
rect 200 59 201 60
rect 201 59 202 60
rect 202 59 203 60
rect 203 59 204 60
rect 204 59 205 60
rect 205 59 206 60
rect 317 59 318 60
rect 318 59 319 60
rect 319 59 320 60
rect 320 59 321 60
rect 321 59 322 60
rect 322 59 323 60
rect 323 59 324 60
rect 394 59 395 60
rect 395 59 396 60
rect 396 59 397 60
rect 397 59 398 60
rect 398 59 399 60
rect 399 59 400 60
rect 400 59 401 60
rect 401 59 402 60
rect 402 59 403 60
rect 403 59 404 60
rect 404 59 405 60
rect 405 59 406 60
rect 182 58 183 59
rect 183 58 184 59
rect 184 58 185 59
rect 185 58 186 59
rect 186 58 187 59
rect 187 58 188 59
rect 188 58 189 59
rect 189 58 190 59
rect 190 58 191 59
rect 191 58 192 59
rect 192 58 193 59
rect 193 58 194 59
rect 194 58 195 59
rect 195 58 196 59
rect 196 58 197 59
rect 197 58 198 59
rect 198 58 199 59
rect 199 58 200 59
rect 200 58 201 59
rect 201 58 202 59
rect 202 58 203 59
rect 203 58 204 59
rect 204 58 205 59
rect 205 58 206 59
rect 206 58 207 59
rect 207 58 208 59
rect 208 58 209 59
rect 311 58 312 59
rect 312 58 313 59
rect 313 58 314 59
rect 314 58 315 59
rect 315 58 316 59
rect 316 58 317 59
rect 317 58 318 59
rect 318 58 319 59
rect 319 58 320 59
rect 320 58 321 59
rect 321 58 322 59
rect 322 58 323 59
rect 323 58 324 59
rect 392 58 393 59
rect 393 58 394 59
rect 394 58 395 59
rect 395 58 396 59
rect 396 58 397 59
rect 397 58 398 59
rect 398 58 399 59
rect 399 58 400 59
rect 400 58 401 59
rect 401 58 402 59
rect 402 58 403 59
rect 403 58 404 59
rect 404 58 405 59
rect 405 58 406 59
rect 186 57 187 58
rect 187 57 188 58
rect 188 57 189 58
rect 189 57 190 58
rect 190 57 191 58
rect 191 57 192 58
rect 192 57 193 58
rect 193 57 194 58
rect 194 57 195 58
rect 195 57 196 58
rect 196 57 197 58
rect 197 57 198 58
rect 198 57 199 58
rect 199 57 200 58
rect 200 57 201 58
rect 201 57 202 58
rect 202 57 203 58
rect 203 57 204 58
rect 204 57 205 58
rect 205 57 206 58
rect 206 57 207 58
rect 207 57 208 58
rect 208 57 209 58
rect 311 57 312 58
rect 312 57 313 58
rect 313 57 314 58
rect 314 57 315 58
rect 315 57 316 58
rect 316 57 317 58
rect 317 57 318 58
rect 318 57 319 58
rect 319 57 320 58
rect 392 57 393 58
rect 393 57 394 58
rect 394 57 395 58
rect 395 57 396 58
rect 396 57 397 58
rect 397 57 398 58
rect 398 57 399 58
rect 399 57 400 58
rect 400 57 401 58
rect 401 57 402 58
rect 186 56 187 57
rect 187 56 188 57
rect 188 56 189 57
rect 189 56 190 57
rect 190 56 191 57
rect 191 56 192 57
rect 192 56 193 57
rect 193 56 194 57
rect 194 56 195 57
rect 195 56 196 57
rect 196 56 197 57
rect 197 56 198 57
rect 198 56 199 57
rect 199 56 200 57
rect 200 56 201 57
rect 201 56 202 57
rect 202 56 203 57
rect 203 56 204 57
rect 204 56 205 57
rect 205 56 206 57
rect 206 56 207 57
rect 207 56 208 57
rect 208 56 209 57
rect 209 56 210 57
rect 210 56 211 57
rect 211 56 212 57
rect 212 56 213 57
rect 213 56 214 57
rect 214 56 215 57
rect 215 56 216 57
rect 216 56 217 57
rect 217 56 218 57
rect 218 56 219 57
rect 219 56 220 57
rect 220 56 221 57
rect 221 56 222 57
rect 223 56 224 57
rect 224 56 225 57
rect 225 56 226 57
rect 300 56 301 57
rect 301 56 302 57
rect 302 56 303 57
rect 304 56 305 57
rect 305 56 306 57
rect 306 56 307 57
rect 307 56 308 57
rect 308 56 309 57
rect 309 56 310 57
rect 310 56 311 57
rect 311 56 312 57
rect 312 56 313 57
rect 313 56 314 57
rect 314 56 315 57
rect 315 56 316 57
rect 316 56 317 57
rect 317 56 318 57
rect 318 56 319 57
rect 319 56 320 57
rect 388 56 389 57
rect 389 56 390 57
rect 390 56 391 57
rect 391 56 392 57
rect 392 56 393 57
rect 393 56 394 57
rect 394 56 395 57
rect 395 56 396 57
rect 396 56 397 57
rect 397 56 398 57
rect 398 56 399 57
rect 399 56 400 57
rect 400 56 401 57
rect 401 56 402 57
rect 188 55 189 56
rect 189 55 190 56
rect 190 55 191 56
rect 191 55 192 56
rect 192 55 193 56
rect 193 55 194 56
rect 194 55 195 56
rect 195 55 196 56
rect 196 55 197 56
rect 197 55 198 56
rect 198 55 199 56
rect 199 55 200 56
rect 200 55 201 56
rect 201 55 202 56
rect 202 55 203 56
rect 203 55 204 56
rect 204 55 205 56
rect 205 55 206 56
rect 206 55 207 56
rect 207 55 208 56
rect 208 55 209 56
rect 209 55 210 56
rect 210 55 211 56
rect 211 55 212 56
rect 212 55 213 56
rect 213 55 214 56
rect 214 55 215 56
rect 215 55 216 56
rect 216 55 217 56
rect 217 55 218 56
rect 218 55 219 56
rect 219 55 220 56
rect 220 55 221 56
rect 221 55 222 56
rect 223 55 224 56
rect 224 55 225 56
rect 225 55 226 56
rect 300 55 301 56
rect 301 55 302 56
rect 302 55 303 56
rect 304 55 305 56
rect 305 55 306 56
rect 306 55 307 56
rect 307 55 308 56
rect 308 55 309 56
rect 309 55 310 56
rect 310 55 311 56
rect 311 55 312 56
rect 312 55 313 56
rect 313 55 314 56
rect 314 55 315 56
rect 315 55 316 56
rect 316 55 317 56
rect 317 55 318 56
rect 388 55 389 56
rect 389 55 390 56
rect 390 55 391 56
rect 391 55 392 56
rect 392 55 393 56
rect 393 55 394 56
rect 394 55 395 56
rect 395 55 396 56
rect 396 55 397 56
rect 397 55 398 56
rect 398 55 399 56
rect 399 55 400 56
rect 188 54 189 55
rect 189 54 190 55
rect 190 54 191 55
rect 191 54 192 55
rect 192 54 193 55
rect 193 54 194 55
rect 194 54 195 55
rect 195 54 196 55
rect 196 54 197 55
rect 197 54 198 55
rect 198 54 199 55
rect 199 54 200 55
rect 200 54 201 55
rect 201 54 202 55
rect 202 54 203 55
rect 203 54 204 55
rect 204 54 205 55
rect 205 54 206 55
rect 206 54 207 55
rect 207 54 208 55
rect 208 54 209 55
rect 209 54 210 55
rect 210 54 211 55
rect 211 54 212 55
rect 212 54 213 55
rect 213 54 214 55
rect 214 54 215 55
rect 215 54 216 55
rect 216 54 217 55
rect 217 54 218 55
rect 218 54 219 55
rect 219 54 220 55
rect 220 54 221 55
rect 221 54 222 55
rect 222 54 223 55
rect 223 54 224 55
rect 224 54 225 55
rect 225 54 226 55
rect 226 54 227 55
rect 227 54 228 55
rect 228 54 229 55
rect 229 54 230 55
rect 230 54 231 55
rect 231 54 232 55
rect 232 54 233 55
rect 233 54 234 55
rect 234 54 235 55
rect 235 54 236 55
rect 236 54 237 55
rect 237 54 238 55
rect 238 54 239 55
rect 240 54 241 55
rect 241 54 242 55
rect 242 54 243 55
rect 244 54 245 55
rect 245 54 246 55
rect 246 54 247 55
rect 248 54 249 55
rect 249 54 250 55
rect 250 54 251 55
rect 279 54 280 55
rect 280 54 281 55
rect 281 54 282 55
rect 285 54 286 55
rect 286 54 287 55
rect 287 54 288 55
rect 289 54 290 55
rect 290 54 291 55
rect 291 54 292 55
rect 292 54 293 55
rect 293 54 294 55
rect 294 54 295 55
rect 295 54 296 55
rect 296 54 297 55
rect 297 54 298 55
rect 298 54 299 55
rect 299 54 300 55
rect 300 54 301 55
rect 301 54 302 55
rect 302 54 303 55
rect 303 54 304 55
rect 304 54 305 55
rect 305 54 306 55
rect 306 54 307 55
rect 307 54 308 55
rect 308 54 309 55
rect 309 54 310 55
rect 310 54 311 55
rect 311 54 312 55
rect 312 54 313 55
rect 313 54 314 55
rect 314 54 315 55
rect 315 54 316 55
rect 316 54 317 55
rect 317 54 318 55
rect 386 54 387 55
rect 387 54 388 55
rect 388 54 389 55
rect 389 54 390 55
rect 390 54 391 55
rect 391 54 392 55
rect 392 54 393 55
rect 393 54 394 55
rect 394 54 395 55
rect 395 54 396 55
rect 396 54 397 55
rect 397 54 398 55
rect 398 54 399 55
rect 399 54 400 55
rect 191 53 192 54
rect 192 53 193 54
rect 193 53 194 54
rect 194 53 195 54
rect 195 53 196 54
rect 196 53 197 54
rect 197 53 198 54
rect 198 53 199 54
rect 199 53 200 54
rect 200 53 201 54
rect 201 53 202 54
rect 202 53 203 54
rect 203 53 204 54
rect 204 53 205 54
rect 205 53 206 54
rect 206 53 207 54
rect 207 53 208 54
rect 208 53 209 54
rect 209 53 210 54
rect 210 53 211 54
rect 211 53 212 54
rect 212 53 213 54
rect 213 53 214 54
rect 214 53 215 54
rect 215 53 216 54
rect 216 53 217 54
rect 217 53 218 54
rect 218 53 219 54
rect 219 53 220 54
rect 220 53 221 54
rect 221 53 222 54
rect 222 53 223 54
rect 223 53 224 54
rect 224 53 225 54
rect 225 53 226 54
rect 226 53 227 54
rect 227 53 228 54
rect 228 53 229 54
rect 229 53 230 54
rect 230 53 231 54
rect 231 53 232 54
rect 232 53 233 54
rect 233 53 234 54
rect 234 53 235 54
rect 235 53 236 54
rect 236 53 237 54
rect 237 53 238 54
rect 238 53 239 54
rect 240 53 241 54
rect 241 53 242 54
rect 242 53 243 54
rect 244 53 245 54
rect 245 53 246 54
rect 246 53 247 54
rect 248 53 249 54
rect 249 53 250 54
rect 250 53 251 54
rect 279 53 280 54
rect 280 53 281 54
rect 281 53 282 54
rect 285 53 286 54
rect 286 53 287 54
rect 287 53 288 54
rect 289 53 290 54
rect 290 53 291 54
rect 291 53 292 54
rect 292 53 293 54
rect 293 53 294 54
rect 294 53 295 54
rect 295 53 296 54
rect 296 53 297 54
rect 297 53 298 54
rect 298 53 299 54
rect 299 53 300 54
rect 300 53 301 54
rect 301 53 302 54
rect 302 53 303 54
rect 303 53 304 54
rect 304 53 305 54
rect 305 53 306 54
rect 306 53 307 54
rect 307 53 308 54
rect 308 53 309 54
rect 309 53 310 54
rect 310 53 311 54
rect 311 53 312 54
rect 312 53 313 54
rect 313 53 314 54
rect 386 53 387 54
rect 387 53 388 54
rect 388 53 389 54
rect 389 53 390 54
rect 390 53 391 54
rect 391 53 392 54
rect 392 53 393 54
rect 393 53 394 54
rect 394 53 395 54
rect 395 53 396 54
rect 396 53 397 54
rect 191 52 192 53
rect 192 52 193 53
rect 193 52 194 53
rect 194 52 195 53
rect 195 52 196 53
rect 196 52 197 53
rect 197 52 198 53
rect 198 52 199 53
rect 199 52 200 53
rect 200 52 201 53
rect 201 52 202 53
rect 202 52 203 53
rect 203 52 204 53
rect 204 52 205 53
rect 205 52 206 53
rect 206 52 207 53
rect 207 52 208 53
rect 208 52 209 53
rect 209 52 210 53
rect 210 52 211 53
rect 211 52 212 53
rect 212 52 213 53
rect 213 52 214 53
rect 214 52 215 53
rect 215 52 216 53
rect 216 52 217 53
rect 217 52 218 53
rect 218 52 219 53
rect 219 52 220 53
rect 220 52 221 53
rect 221 52 222 53
rect 222 52 223 53
rect 223 52 224 53
rect 224 52 225 53
rect 225 52 226 53
rect 226 52 227 53
rect 227 52 228 53
rect 228 52 229 53
rect 229 52 230 53
rect 230 52 231 53
rect 231 52 232 53
rect 232 52 233 53
rect 233 52 234 53
rect 234 52 235 53
rect 235 52 236 53
rect 236 52 237 53
rect 237 52 238 53
rect 238 52 239 53
rect 239 52 240 53
rect 240 52 241 53
rect 241 52 242 53
rect 242 52 243 53
rect 243 52 244 53
rect 244 52 245 53
rect 245 52 246 53
rect 246 52 247 53
rect 247 52 248 53
rect 248 52 249 53
rect 249 52 250 53
rect 250 52 251 53
rect 251 52 252 53
rect 252 52 253 53
rect 253 52 254 53
rect 254 52 255 53
rect 255 52 256 53
rect 256 52 257 53
rect 257 52 258 53
rect 258 52 259 53
rect 259 52 260 53
rect 260 52 261 53
rect 261 52 262 53
rect 262 52 263 53
rect 263 52 264 53
rect 264 52 265 53
rect 265 52 266 53
rect 266 52 267 53
rect 267 52 268 53
rect 268 52 269 53
rect 269 52 270 53
rect 270 52 271 53
rect 271 52 272 53
rect 272 52 273 53
rect 273 52 274 53
rect 274 52 275 53
rect 275 52 276 53
rect 276 52 277 53
rect 277 52 278 53
rect 278 52 279 53
rect 279 52 280 53
rect 280 52 281 53
rect 281 52 282 53
rect 282 52 283 53
rect 283 52 284 53
rect 284 52 285 53
rect 285 52 286 53
rect 286 52 287 53
rect 287 52 288 53
rect 288 52 289 53
rect 289 52 290 53
rect 290 52 291 53
rect 291 52 292 53
rect 292 52 293 53
rect 293 52 294 53
rect 294 52 295 53
rect 295 52 296 53
rect 296 52 297 53
rect 297 52 298 53
rect 298 52 299 53
rect 299 52 300 53
rect 300 52 301 53
rect 301 52 302 53
rect 302 52 303 53
rect 303 52 304 53
rect 304 52 305 53
rect 305 52 306 53
rect 306 52 307 53
rect 307 52 308 53
rect 308 52 309 53
rect 309 52 310 53
rect 310 52 311 53
rect 311 52 312 53
rect 312 52 313 53
rect 313 52 314 53
rect 383 52 384 53
rect 384 52 385 53
rect 385 52 386 53
rect 386 52 387 53
rect 387 52 388 53
rect 388 52 389 53
rect 389 52 390 53
rect 390 52 391 53
rect 391 52 392 53
rect 392 52 393 53
rect 393 52 394 53
rect 394 52 395 53
rect 395 52 396 53
rect 396 52 397 53
rect 195 51 196 52
rect 196 51 197 52
rect 197 51 198 52
rect 198 51 199 52
rect 199 51 200 52
rect 200 51 201 52
rect 201 51 202 52
rect 202 51 203 52
rect 203 51 204 52
rect 204 51 205 52
rect 205 51 206 52
rect 206 51 207 52
rect 207 51 208 52
rect 208 51 209 52
rect 209 51 210 52
rect 210 51 211 52
rect 211 51 212 52
rect 212 51 213 52
rect 213 51 214 52
rect 214 51 215 52
rect 215 51 216 52
rect 216 51 217 52
rect 217 51 218 52
rect 218 51 219 52
rect 219 51 220 52
rect 220 51 221 52
rect 221 51 222 52
rect 222 51 223 52
rect 223 51 224 52
rect 224 51 225 52
rect 225 51 226 52
rect 226 51 227 52
rect 227 51 228 52
rect 228 51 229 52
rect 229 51 230 52
rect 230 51 231 52
rect 231 51 232 52
rect 232 51 233 52
rect 233 51 234 52
rect 234 51 235 52
rect 235 51 236 52
rect 236 51 237 52
rect 237 51 238 52
rect 238 51 239 52
rect 239 51 240 52
rect 240 51 241 52
rect 241 51 242 52
rect 242 51 243 52
rect 243 51 244 52
rect 244 51 245 52
rect 245 51 246 52
rect 246 51 247 52
rect 247 51 248 52
rect 248 51 249 52
rect 249 51 250 52
rect 250 51 251 52
rect 251 51 252 52
rect 252 51 253 52
rect 253 51 254 52
rect 254 51 255 52
rect 255 51 256 52
rect 256 51 257 52
rect 257 51 258 52
rect 258 51 259 52
rect 259 51 260 52
rect 260 51 261 52
rect 261 51 262 52
rect 262 51 263 52
rect 263 51 264 52
rect 264 51 265 52
rect 265 51 266 52
rect 266 51 267 52
rect 267 51 268 52
rect 268 51 269 52
rect 269 51 270 52
rect 270 51 271 52
rect 271 51 272 52
rect 272 51 273 52
rect 273 51 274 52
rect 274 51 275 52
rect 275 51 276 52
rect 276 51 277 52
rect 277 51 278 52
rect 278 51 279 52
rect 279 51 280 52
rect 280 51 281 52
rect 281 51 282 52
rect 282 51 283 52
rect 283 51 284 52
rect 284 51 285 52
rect 285 51 286 52
rect 286 51 287 52
rect 287 51 288 52
rect 288 51 289 52
rect 289 51 290 52
rect 290 51 291 52
rect 291 51 292 52
rect 292 51 293 52
rect 293 51 294 52
rect 294 51 295 52
rect 295 51 296 52
rect 296 51 297 52
rect 297 51 298 52
rect 298 51 299 52
rect 299 51 300 52
rect 300 51 301 52
rect 301 51 302 52
rect 302 51 303 52
rect 303 51 304 52
rect 304 51 305 52
rect 305 51 306 52
rect 306 51 307 52
rect 307 51 308 52
rect 308 51 309 52
rect 309 51 310 52
rect 310 51 311 52
rect 311 51 312 52
rect 383 51 384 52
rect 384 51 385 52
rect 385 51 386 52
rect 386 51 387 52
rect 387 51 388 52
rect 388 51 389 52
rect 389 51 390 52
rect 390 51 391 52
rect 391 51 392 52
rect 392 51 393 52
rect 393 51 394 52
rect 394 51 395 52
rect 195 50 196 51
rect 196 50 197 51
rect 197 50 198 51
rect 198 50 199 51
rect 199 50 200 51
rect 200 50 201 51
rect 201 50 202 51
rect 202 50 203 51
rect 203 50 204 51
rect 204 50 205 51
rect 205 50 206 51
rect 206 50 207 51
rect 207 50 208 51
rect 208 50 209 51
rect 209 50 210 51
rect 210 50 211 51
rect 211 50 212 51
rect 212 50 213 51
rect 213 50 214 51
rect 214 50 215 51
rect 215 50 216 51
rect 216 50 217 51
rect 217 50 218 51
rect 218 50 219 51
rect 219 50 220 51
rect 220 50 221 51
rect 221 50 222 51
rect 222 50 223 51
rect 223 50 224 51
rect 224 50 225 51
rect 225 50 226 51
rect 226 50 227 51
rect 227 50 228 51
rect 228 50 229 51
rect 229 50 230 51
rect 230 50 231 51
rect 231 50 232 51
rect 232 50 233 51
rect 233 50 234 51
rect 234 50 235 51
rect 235 50 236 51
rect 236 50 237 51
rect 237 50 238 51
rect 238 50 239 51
rect 239 50 240 51
rect 240 50 241 51
rect 241 50 242 51
rect 242 50 243 51
rect 243 50 244 51
rect 244 50 245 51
rect 245 50 246 51
rect 246 50 247 51
rect 247 50 248 51
rect 248 50 249 51
rect 249 50 250 51
rect 250 50 251 51
rect 251 50 252 51
rect 252 50 253 51
rect 253 50 254 51
rect 254 50 255 51
rect 255 50 256 51
rect 256 50 257 51
rect 257 50 258 51
rect 258 50 259 51
rect 259 50 260 51
rect 260 50 261 51
rect 261 50 262 51
rect 262 50 263 51
rect 263 50 264 51
rect 264 50 265 51
rect 265 50 266 51
rect 266 50 267 51
rect 267 50 268 51
rect 268 50 269 51
rect 269 50 270 51
rect 270 50 271 51
rect 271 50 272 51
rect 272 50 273 51
rect 273 50 274 51
rect 274 50 275 51
rect 275 50 276 51
rect 276 50 277 51
rect 277 50 278 51
rect 278 50 279 51
rect 279 50 280 51
rect 280 50 281 51
rect 281 50 282 51
rect 282 50 283 51
rect 283 50 284 51
rect 284 50 285 51
rect 285 50 286 51
rect 286 50 287 51
rect 287 50 288 51
rect 288 50 289 51
rect 289 50 290 51
rect 290 50 291 51
rect 291 50 292 51
rect 292 50 293 51
rect 293 50 294 51
rect 294 50 295 51
rect 295 50 296 51
rect 296 50 297 51
rect 297 50 298 51
rect 298 50 299 51
rect 299 50 300 51
rect 300 50 301 51
rect 301 50 302 51
rect 302 50 303 51
rect 303 50 304 51
rect 304 50 305 51
rect 305 50 306 51
rect 306 50 307 51
rect 307 50 308 51
rect 308 50 309 51
rect 309 50 310 51
rect 310 50 311 51
rect 311 50 312 51
rect 381 50 382 51
rect 382 50 383 51
rect 383 50 384 51
rect 384 50 385 51
rect 385 50 386 51
rect 386 50 387 51
rect 387 50 388 51
rect 388 50 389 51
rect 389 50 390 51
rect 390 50 391 51
rect 391 50 392 51
rect 392 50 393 51
rect 393 50 394 51
rect 394 50 395 51
rect 199 49 200 50
rect 200 49 201 50
rect 201 49 202 50
rect 202 49 203 50
rect 203 49 204 50
rect 204 49 205 50
rect 205 49 206 50
rect 206 49 207 50
rect 207 49 208 50
rect 208 49 209 50
rect 209 49 210 50
rect 210 49 211 50
rect 211 49 212 50
rect 212 49 213 50
rect 213 49 214 50
rect 214 49 215 50
rect 215 49 216 50
rect 216 49 217 50
rect 217 49 218 50
rect 218 49 219 50
rect 219 49 220 50
rect 220 49 221 50
rect 221 49 222 50
rect 222 49 223 50
rect 223 49 224 50
rect 224 49 225 50
rect 225 49 226 50
rect 226 49 227 50
rect 227 49 228 50
rect 228 49 229 50
rect 229 49 230 50
rect 230 49 231 50
rect 231 49 232 50
rect 232 49 233 50
rect 233 49 234 50
rect 234 49 235 50
rect 235 49 236 50
rect 236 49 237 50
rect 237 49 238 50
rect 238 49 239 50
rect 239 49 240 50
rect 240 49 241 50
rect 241 49 242 50
rect 242 49 243 50
rect 243 49 244 50
rect 244 49 245 50
rect 245 49 246 50
rect 246 49 247 50
rect 247 49 248 50
rect 248 49 249 50
rect 249 49 250 50
rect 250 49 251 50
rect 251 49 252 50
rect 252 49 253 50
rect 253 49 254 50
rect 254 49 255 50
rect 255 49 256 50
rect 256 49 257 50
rect 257 49 258 50
rect 258 49 259 50
rect 259 49 260 50
rect 260 49 261 50
rect 261 49 262 50
rect 262 49 263 50
rect 263 49 264 50
rect 264 49 265 50
rect 265 49 266 50
rect 266 49 267 50
rect 267 49 268 50
rect 268 49 269 50
rect 269 49 270 50
rect 270 49 271 50
rect 271 49 272 50
rect 272 49 273 50
rect 273 49 274 50
rect 274 49 275 50
rect 275 49 276 50
rect 276 49 277 50
rect 277 49 278 50
rect 278 49 279 50
rect 279 49 280 50
rect 280 49 281 50
rect 281 49 282 50
rect 282 49 283 50
rect 283 49 284 50
rect 284 49 285 50
rect 285 49 286 50
rect 286 49 287 50
rect 287 49 288 50
rect 288 49 289 50
rect 289 49 290 50
rect 290 49 291 50
rect 291 49 292 50
rect 292 49 293 50
rect 293 49 294 50
rect 294 49 295 50
rect 295 49 296 50
rect 296 49 297 50
rect 297 49 298 50
rect 298 49 299 50
rect 299 49 300 50
rect 300 49 301 50
rect 301 49 302 50
rect 302 49 303 50
rect 303 49 304 50
rect 304 49 305 50
rect 305 49 306 50
rect 306 49 307 50
rect 307 49 308 50
rect 308 49 309 50
rect 309 49 310 50
rect 381 49 382 50
rect 382 49 383 50
rect 383 49 384 50
rect 384 49 385 50
rect 385 49 386 50
rect 386 49 387 50
rect 387 49 388 50
rect 388 49 389 50
rect 389 49 390 50
rect 390 49 391 50
rect 199 48 200 49
rect 200 48 201 49
rect 201 48 202 49
rect 202 48 203 49
rect 203 48 204 49
rect 204 48 205 49
rect 205 48 206 49
rect 206 48 207 49
rect 207 48 208 49
rect 208 48 209 49
rect 209 48 210 49
rect 210 48 211 49
rect 211 48 212 49
rect 212 48 213 49
rect 213 48 214 49
rect 214 48 215 49
rect 215 48 216 49
rect 216 48 217 49
rect 217 48 218 49
rect 218 48 219 49
rect 219 48 220 49
rect 220 48 221 49
rect 221 48 222 49
rect 222 48 223 49
rect 223 48 224 49
rect 224 48 225 49
rect 225 48 226 49
rect 226 48 227 49
rect 227 48 228 49
rect 228 48 229 49
rect 229 48 230 49
rect 230 48 231 49
rect 231 48 232 49
rect 232 48 233 49
rect 233 48 234 49
rect 234 48 235 49
rect 235 48 236 49
rect 236 48 237 49
rect 237 48 238 49
rect 238 48 239 49
rect 239 48 240 49
rect 240 48 241 49
rect 241 48 242 49
rect 242 48 243 49
rect 243 48 244 49
rect 244 48 245 49
rect 245 48 246 49
rect 246 48 247 49
rect 247 48 248 49
rect 248 48 249 49
rect 249 48 250 49
rect 250 48 251 49
rect 251 48 252 49
rect 252 48 253 49
rect 253 48 254 49
rect 254 48 255 49
rect 255 48 256 49
rect 256 48 257 49
rect 257 48 258 49
rect 258 48 259 49
rect 259 48 260 49
rect 260 48 261 49
rect 261 48 262 49
rect 262 48 263 49
rect 263 48 264 49
rect 264 48 265 49
rect 265 48 266 49
rect 266 48 267 49
rect 267 48 268 49
rect 268 48 269 49
rect 269 48 270 49
rect 270 48 271 49
rect 271 48 272 49
rect 272 48 273 49
rect 273 48 274 49
rect 274 48 275 49
rect 275 48 276 49
rect 276 48 277 49
rect 277 48 278 49
rect 278 48 279 49
rect 279 48 280 49
rect 280 48 281 49
rect 281 48 282 49
rect 282 48 283 49
rect 283 48 284 49
rect 284 48 285 49
rect 285 48 286 49
rect 286 48 287 49
rect 287 48 288 49
rect 288 48 289 49
rect 289 48 290 49
rect 290 48 291 49
rect 291 48 292 49
rect 292 48 293 49
rect 293 48 294 49
rect 294 48 295 49
rect 295 48 296 49
rect 296 48 297 49
rect 297 48 298 49
rect 298 48 299 49
rect 299 48 300 49
rect 300 48 301 49
rect 301 48 302 49
rect 302 48 303 49
rect 303 48 304 49
rect 304 48 305 49
rect 305 48 306 49
rect 306 48 307 49
rect 307 48 308 49
rect 308 48 309 49
rect 309 48 310 49
rect 310 48 311 49
rect 311 48 312 49
rect 377 48 378 49
rect 378 48 379 49
rect 379 48 380 49
rect 380 48 381 49
rect 381 48 382 49
rect 382 48 383 49
rect 383 48 384 49
rect 384 48 385 49
rect 385 48 386 49
rect 386 48 387 49
rect 387 48 388 49
rect 388 48 389 49
rect 389 48 390 49
rect 390 48 391 49
rect 203 47 204 48
rect 204 47 205 48
rect 205 47 206 48
rect 206 47 207 48
rect 207 47 208 48
rect 208 47 209 48
rect 209 47 210 48
rect 210 47 211 48
rect 211 47 212 48
rect 212 47 213 48
rect 213 47 214 48
rect 214 47 215 48
rect 215 47 216 48
rect 216 47 217 48
rect 217 47 218 48
rect 218 47 219 48
rect 219 47 220 48
rect 220 47 221 48
rect 221 47 222 48
rect 222 47 223 48
rect 223 47 224 48
rect 224 47 225 48
rect 225 47 226 48
rect 226 47 227 48
rect 227 47 228 48
rect 228 47 229 48
rect 229 47 230 48
rect 230 47 231 48
rect 231 47 232 48
rect 232 47 233 48
rect 233 47 234 48
rect 234 47 235 48
rect 235 47 236 48
rect 236 47 237 48
rect 237 47 238 48
rect 238 47 239 48
rect 239 47 240 48
rect 240 47 241 48
rect 241 47 242 48
rect 242 47 243 48
rect 243 47 244 48
rect 244 47 245 48
rect 245 47 246 48
rect 246 47 247 48
rect 247 47 248 48
rect 248 47 249 48
rect 249 47 250 48
rect 250 47 251 48
rect 251 47 252 48
rect 252 47 253 48
rect 253 47 254 48
rect 254 47 255 48
rect 255 47 256 48
rect 256 47 257 48
rect 257 47 258 48
rect 258 47 259 48
rect 259 47 260 48
rect 260 47 261 48
rect 261 47 262 48
rect 262 47 263 48
rect 263 47 264 48
rect 264 47 265 48
rect 265 47 266 48
rect 266 47 267 48
rect 267 47 268 48
rect 268 47 269 48
rect 269 47 270 48
rect 270 47 271 48
rect 271 47 272 48
rect 272 47 273 48
rect 273 47 274 48
rect 274 47 275 48
rect 275 47 276 48
rect 276 47 277 48
rect 277 47 278 48
rect 278 47 279 48
rect 279 47 280 48
rect 280 47 281 48
rect 281 47 282 48
rect 282 47 283 48
rect 283 47 284 48
rect 284 47 285 48
rect 285 47 286 48
rect 286 47 287 48
rect 287 47 288 48
rect 288 47 289 48
rect 289 47 290 48
rect 290 47 291 48
rect 291 47 292 48
rect 292 47 293 48
rect 293 47 294 48
rect 294 47 295 48
rect 295 47 296 48
rect 296 47 297 48
rect 297 47 298 48
rect 298 47 299 48
rect 299 47 300 48
rect 300 47 301 48
rect 301 47 302 48
rect 302 47 303 48
rect 303 47 304 48
rect 304 47 305 48
rect 305 47 306 48
rect 306 47 307 48
rect 307 47 308 48
rect 308 47 309 48
rect 309 47 310 48
rect 310 47 311 48
rect 311 47 312 48
rect 377 47 378 48
rect 378 47 379 48
rect 379 47 380 48
rect 380 47 381 48
rect 381 47 382 48
rect 382 47 383 48
rect 383 47 384 48
rect 384 47 385 48
rect 385 47 386 48
rect 386 47 387 48
rect 387 47 388 48
rect 388 47 389 48
rect 203 46 204 47
rect 204 46 205 47
rect 205 46 206 47
rect 206 46 207 47
rect 207 46 208 47
rect 208 46 209 47
rect 209 46 210 47
rect 210 46 211 47
rect 211 46 212 47
rect 212 46 213 47
rect 213 46 214 47
rect 214 46 215 47
rect 215 46 216 47
rect 216 46 217 47
rect 217 46 218 47
rect 218 46 219 47
rect 219 46 220 47
rect 220 46 221 47
rect 221 46 222 47
rect 222 46 223 47
rect 223 46 224 47
rect 224 46 225 47
rect 225 46 226 47
rect 226 46 227 47
rect 227 46 228 47
rect 228 46 229 47
rect 229 46 230 47
rect 230 46 231 47
rect 231 46 232 47
rect 232 46 233 47
rect 233 46 234 47
rect 234 46 235 47
rect 235 46 236 47
rect 236 46 237 47
rect 237 46 238 47
rect 238 46 239 47
rect 239 46 240 47
rect 240 46 241 47
rect 241 46 242 47
rect 242 46 243 47
rect 243 46 244 47
rect 244 46 245 47
rect 245 46 246 47
rect 246 46 247 47
rect 247 46 248 47
rect 248 46 249 47
rect 249 46 250 47
rect 250 46 251 47
rect 251 46 252 47
rect 252 46 253 47
rect 253 46 254 47
rect 254 46 255 47
rect 255 46 256 47
rect 256 46 257 47
rect 257 46 258 47
rect 258 46 259 47
rect 259 46 260 47
rect 260 46 261 47
rect 261 46 262 47
rect 262 46 263 47
rect 263 46 264 47
rect 264 46 265 47
rect 265 46 266 47
rect 266 46 267 47
rect 267 46 268 47
rect 268 46 269 47
rect 269 46 270 47
rect 270 46 271 47
rect 271 46 272 47
rect 272 46 273 47
rect 273 46 274 47
rect 274 46 275 47
rect 275 46 276 47
rect 276 46 277 47
rect 277 46 278 47
rect 278 46 279 47
rect 279 46 280 47
rect 280 46 281 47
rect 281 46 282 47
rect 282 46 283 47
rect 283 46 284 47
rect 284 46 285 47
rect 285 46 286 47
rect 286 46 287 47
rect 287 46 288 47
rect 288 46 289 47
rect 289 46 290 47
rect 290 46 291 47
rect 291 46 292 47
rect 292 46 293 47
rect 293 46 294 47
rect 294 46 295 47
rect 295 46 296 47
rect 296 46 297 47
rect 297 46 298 47
rect 298 46 299 47
rect 299 46 300 47
rect 300 46 301 47
rect 301 46 302 47
rect 302 46 303 47
rect 303 46 304 47
rect 304 46 305 47
rect 305 46 306 47
rect 306 46 307 47
rect 307 46 308 47
rect 308 46 309 47
rect 309 46 310 47
rect 310 46 311 47
rect 311 46 312 47
rect 312 46 313 47
rect 313 46 314 47
rect 314 46 315 47
rect 315 46 316 47
rect 373 46 374 47
rect 374 46 375 47
rect 375 46 376 47
rect 376 46 377 47
rect 377 46 378 47
rect 378 46 379 47
rect 379 46 380 47
rect 380 46 381 47
rect 381 46 382 47
rect 382 46 383 47
rect 383 46 384 47
rect 384 46 385 47
rect 385 46 386 47
rect 386 46 387 47
rect 387 46 388 47
rect 388 46 389 47
rect 206 45 207 46
rect 207 45 208 46
rect 208 45 209 46
rect 209 45 210 46
rect 210 45 211 46
rect 211 45 212 46
rect 212 45 213 46
rect 213 45 214 46
rect 214 45 215 46
rect 215 45 216 46
rect 216 45 217 46
rect 217 45 218 46
rect 218 45 219 46
rect 219 45 220 46
rect 220 45 221 46
rect 221 45 222 46
rect 222 45 223 46
rect 223 45 224 46
rect 224 45 225 46
rect 225 45 226 46
rect 226 45 227 46
rect 227 45 228 46
rect 228 45 229 46
rect 229 45 230 46
rect 230 45 231 46
rect 231 45 232 46
rect 232 45 233 46
rect 233 45 234 46
rect 234 45 235 46
rect 235 45 236 46
rect 236 45 237 46
rect 237 45 238 46
rect 238 45 239 46
rect 239 45 240 46
rect 240 45 241 46
rect 241 45 242 46
rect 242 45 243 46
rect 243 45 244 46
rect 244 45 245 46
rect 245 45 246 46
rect 246 45 247 46
rect 247 45 248 46
rect 248 45 249 46
rect 249 45 250 46
rect 250 45 251 46
rect 251 45 252 46
rect 252 45 253 46
rect 253 45 254 46
rect 254 45 255 46
rect 255 45 256 46
rect 256 45 257 46
rect 257 45 258 46
rect 258 45 259 46
rect 259 45 260 46
rect 260 45 261 46
rect 261 45 262 46
rect 262 45 263 46
rect 263 45 264 46
rect 264 45 265 46
rect 265 45 266 46
rect 266 45 267 46
rect 267 45 268 46
rect 268 45 269 46
rect 269 45 270 46
rect 270 45 271 46
rect 271 45 272 46
rect 272 45 273 46
rect 273 45 274 46
rect 274 45 275 46
rect 275 45 276 46
rect 276 45 277 46
rect 277 45 278 46
rect 278 45 279 46
rect 279 45 280 46
rect 280 45 281 46
rect 281 45 282 46
rect 282 45 283 46
rect 283 45 284 46
rect 284 45 285 46
rect 285 45 286 46
rect 286 45 287 46
rect 287 45 288 46
rect 288 45 289 46
rect 289 45 290 46
rect 290 45 291 46
rect 291 45 292 46
rect 292 45 293 46
rect 293 45 294 46
rect 294 45 295 46
rect 295 45 296 46
rect 296 45 297 46
rect 297 45 298 46
rect 298 45 299 46
rect 299 45 300 46
rect 300 45 301 46
rect 301 45 302 46
rect 302 45 303 46
rect 303 45 304 46
rect 304 45 305 46
rect 305 45 306 46
rect 306 45 307 46
rect 307 45 308 46
rect 308 45 309 46
rect 309 45 310 46
rect 310 45 311 46
rect 311 45 312 46
rect 312 45 313 46
rect 313 45 314 46
rect 314 45 315 46
rect 315 45 316 46
rect 373 45 374 46
rect 374 45 375 46
rect 375 45 376 46
rect 376 45 377 46
rect 377 45 378 46
rect 378 45 379 46
rect 379 45 380 46
rect 380 45 381 46
rect 381 45 382 46
rect 382 45 383 46
rect 383 45 384 46
rect 384 45 385 46
rect 206 44 207 45
rect 207 44 208 45
rect 208 44 209 45
rect 209 44 210 45
rect 210 44 211 45
rect 211 44 212 45
rect 212 44 213 45
rect 213 44 214 45
rect 214 44 215 45
rect 215 44 216 45
rect 216 44 217 45
rect 217 44 218 45
rect 218 44 219 45
rect 219 44 220 45
rect 220 44 221 45
rect 221 44 222 45
rect 222 44 223 45
rect 223 44 224 45
rect 224 44 225 45
rect 225 44 226 45
rect 226 44 227 45
rect 227 44 228 45
rect 228 44 229 45
rect 229 44 230 45
rect 230 44 231 45
rect 231 44 232 45
rect 232 44 233 45
rect 233 44 234 45
rect 234 44 235 45
rect 235 44 236 45
rect 236 44 237 45
rect 237 44 238 45
rect 238 44 239 45
rect 239 44 240 45
rect 240 44 241 45
rect 241 44 242 45
rect 242 44 243 45
rect 243 44 244 45
rect 244 44 245 45
rect 245 44 246 45
rect 246 44 247 45
rect 247 44 248 45
rect 248 44 249 45
rect 249 44 250 45
rect 250 44 251 45
rect 251 44 252 45
rect 252 44 253 45
rect 253 44 254 45
rect 254 44 255 45
rect 255 44 256 45
rect 256 44 257 45
rect 257 44 258 45
rect 258 44 259 45
rect 259 44 260 45
rect 260 44 261 45
rect 261 44 262 45
rect 262 44 263 45
rect 263 44 264 45
rect 264 44 265 45
rect 265 44 266 45
rect 266 44 267 45
rect 267 44 268 45
rect 268 44 269 45
rect 269 44 270 45
rect 270 44 271 45
rect 271 44 272 45
rect 272 44 273 45
rect 273 44 274 45
rect 274 44 275 45
rect 275 44 276 45
rect 276 44 277 45
rect 277 44 278 45
rect 278 44 279 45
rect 279 44 280 45
rect 280 44 281 45
rect 281 44 282 45
rect 282 44 283 45
rect 283 44 284 45
rect 284 44 285 45
rect 285 44 286 45
rect 286 44 287 45
rect 287 44 288 45
rect 288 44 289 45
rect 289 44 290 45
rect 290 44 291 45
rect 291 44 292 45
rect 292 44 293 45
rect 293 44 294 45
rect 294 44 295 45
rect 295 44 296 45
rect 296 44 297 45
rect 297 44 298 45
rect 298 44 299 45
rect 299 44 300 45
rect 300 44 301 45
rect 301 44 302 45
rect 302 44 303 45
rect 303 44 304 45
rect 304 44 305 45
rect 305 44 306 45
rect 306 44 307 45
rect 307 44 308 45
rect 308 44 309 45
rect 309 44 310 45
rect 310 44 311 45
rect 311 44 312 45
rect 312 44 313 45
rect 313 44 314 45
rect 314 44 315 45
rect 315 44 316 45
rect 316 44 317 45
rect 317 44 318 45
rect 318 44 319 45
rect 319 44 320 45
rect 369 44 370 45
rect 370 44 371 45
rect 371 44 372 45
rect 372 44 373 45
rect 373 44 374 45
rect 374 44 375 45
rect 375 44 376 45
rect 376 44 377 45
rect 377 44 378 45
rect 378 44 379 45
rect 379 44 380 45
rect 380 44 381 45
rect 381 44 382 45
rect 382 44 383 45
rect 383 44 384 45
rect 384 44 385 45
rect 210 43 211 44
rect 211 43 212 44
rect 212 43 213 44
rect 213 43 214 44
rect 214 43 215 44
rect 215 43 216 44
rect 216 43 217 44
rect 217 43 218 44
rect 218 43 219 44
rect 219 43 220 44
rect 220 43 221 44
rect 221 43 222 44
rect 222 43 223 44
rect 223 43 224 44
rect 224 43 225 44
rect 225 43 226 44
rect 226 43 227 44
rect 227 43 228 44
rect 228 43 229 44
rect 229 43 230 44
rect 231 43 232 44
rect 232 43 233 44
rect 233 43 234 44
rect 235 43 236 44
rect 236 43 237 44
rect 238 43 239 44
rect 239 43 240 44
rect 240 43 241 44
rect 242 43 243 44
rect 243 43 244 44
rect 244 43 245 44
rect 246 43 247 44
rect 247 43 248 44
rect 248 43 249 44
rect 249 43 250 44
rect 250 43 251 44
rect 251 43 252 44
rect 252 43 253 44
rect 253 43 254 44
rect 254 43 255 44
rect 255 43 256 44
rect 256 43 257 44
rect 257 43 258 44
rect 258 43 259 44
rect 259 43 260 44
rect 260 43 261 44
rect 261 43 262 44
rect 262 43 263 44
rect 263 43 264 44
rect 264 43 265 44
rect 265 43 266 44
rect 266 43 267 44
rect 267 43 268 44
rect 268 43 269 44
rect 269 43 270 44
rect 270 43 271 44
rect 271 43 272 44
rect 272 43 273 44
rect 273 43 274 44
rect 274 43 275 44
rect 275 43 276 44
rect 276 43 277 44
rect 277 43 278 44
rect 278 43 279 44
rect 279 43 280 44
rect 280 43 281 44
rect 281 43 282 44
rect 282 43 283 44
rect 283 43 284 44
rect 284 43 285 44
rect 285 43 286 44
rect 286 43 287 44
rect 287 43 288 44
rect 288 43 289 44
rect 289 43 290 44
rect 290 43 291 44
rect 291 43 292 44
rect 292 43 293 44
rect 293 43 294 44
rect 294 43 295 44
rect 295 43 296 44
rect 296 43 297 44
rect 297 43 298 44
rect 298 43 299 44
rect 299 43 300 44
rect 300 43 301 44
rect 301 43 302 44
rect 302 43 303 44
rect 303 43 304 44
rect 304 43 305 44
rect 305 43 306 44
rect 306 43 307 44
rect 307 43 308 44
rect 308 43 309 44
rect 309 43 310 44
rect 310 43 311 44
rect 311 43 312 44
rect 312 43 313 44
rect 313 43 314 44
rect 314 43 315 44
rect 315 43 316 44
rect 316 43 317 44
rect 317 43 318 44
rect 318 43 319 44
rect 319 43 320 44
rect 369 43 370 44
rect 370 43 371 44
rect 371 43 372 44
rect 372 43 373 44
rect 373 43 374 44
rect 374 43 375 44
rect 375 43 376 44
rect 376 43 377 44
rect 377 43 378 44
rect 378 43 379 44
rect 379 43 380 44
rect 380 43 381 44
rect 381 43 382 44
rect 382 43 383 44
rect 383 43 384 44
rect 210 42 211 43
rect 211 42 212 43
rect 212 42 213 43
rect 213 42 214 43
rect 214 42 215 43
rect 215 42 216 43
rect 216 42 217 43
rect 217 42 218 43
rect 218 42 219 43
rect 219 42 220 43
rect 220 42 221 43
rect 221 42 222 43
rect 222 42 223 43
rect 223 42 224 43
rect 224 42 225 43
rect 225 42 226 43
rect 226 42 227 43
rect 227 42 228 43
rect 228 42 229 43
rect 229 42 230 43
rect 231 42 232 43
rect 232 42 233 43
rect 233 42 234 43
rect 235 42 236 43
rect 236 42 237 43
rect 238 42 239 43
rect 239 42 240 43
rect 240 42 241 43
rect 242 42 243 43
rect 243 42 244 43
rect 244 42 245 43
rect 246 42 247 43
rect 247 42 248 43
rect 248 42 249 43
rect 249 42 250 43
rect 250 42 251 43
rect 251 42 252 43
rect 252 42 253 43
rect 253 42 254 43
rect 254 42 255 43
rect 255 42 256 43
rect 256 42 257 43
rect 257 42 258 43
rect 258 42 259 43
rect 259 42 260 43
rect 260 42 261 43
rect 261 42 262 43
rect 262 42 263 43
rect 263 42 264 43
rect 264 42 265 43
rect 265 42 266 43
rect 266 42 267 43
rect 267 42 268 43
rect 268 42 269 43
rect 269 42 270 43
rect 270 42 271 43
rect 271 42 272 43
rect 272 42 273 43
rect 273 42 274 43
rect 274 42 275 43
rect 275 42 276 43
rect 276 42 277 43
rect 277 42 278 43
rect 278 42 279 43
rect 279 42 280 43
rect 280 42 281 43
rect 281 42 282 43
rect 282 42 283 43
rect 283 42 284 43
rect 284 42 285 43
rect 285 42 286 43
rect 286 42 287 43
rect 287 42 288 43
rect 288 42 289 43
rect 289 42 290 43
rect 290 42 291 43
rect 291 42 292 43
rect 292 42 293 43
rect 293 42 294 43
rect 294 42 295 43
rect 295 42 296 43
rect 296 42 297 43
rect 297 42 298 43
rect 298 42 299 43
rect 299 42 300 43
rect 300 42 301 43
rect 301 42 302 43
rect 302 42 303 43
rect 303 42 304 43
rect 304 42 305 43
rect 305 42 306 43
rect 306 42 307 43
rect 307 42 308 43
rect 308 42 309 43
rect 309 42 310 43
rect 310 42 311 43
rect 311 42 312 43
rect 312 42 313 43
rect 313 42 314 43
rect 314 42 315 43
rect 315 42 316 43
rect 316 42 317 43
rect 317 42 318 43
rect 318 42 319 43
rect 319 42 320 43
rect 320 42 321 43
rect 321 42 322 43
rect 322 42 323 43
rect 323 42 324 43
rect 366 42 367 43
rect 367 42 368 43
rect 368 42 369 43
rect 369 42 370 43
rect 370 42 371 43
rect 371 42 372 43
rect 372 42 373 43
rect 373 42 374 43
rect 374 42 375 43
rect 375 42 376 43
rect 376 42 377 43
rect 377 42 378 43
rect 378 42 379 43
rect 379 42 380 43
rect 380 42 381 43
rect 381 42 382 43
rect 382 42 383 43
rect 383 42 384 43
rect 214 41 215 42
rect 215 41 216 42
rect 216 41 217 42
rect 255 41 256 42
rect 256 41 257 42
rect 257 41 258 42
rect 258 41 259 42
rect 259 41 260 42
rect 260 41 261 42
rect 261 41 262 42
rect 262 41 263 42
rect 263 41 264 42
rect 264 41 265 42
rect 265 41 266 42
rect 266 41 267 42
rect 267 41 268 42
rect 268 41 269 42
rect 269 41 270 42
rect 270 41 271 42
rect 271 41 272 42
rect 272 41 273 42
rect 273 41 274 42
rect 274 41 275 42
rect 275 41 276 42
rect 276 41 277 42
rect 277 41 278 42
rect 278 41 279 42
rect 279 41 280 42
rect 280 41 281 42
rect 281 41 282 42
rect 282 41 283 42
rect 283 41 284 42
rect 284 41 285 42
rect 285 41 286 42
rect 286 41 287 42
rect 287 41 288 42
rect 288 41 289 42
rect 289 41 290 42
rect 290 41 291 42
rect 291 41 292 42
rect 292 41 293 42
rect 293 41 294 42
rect 294 41 295 42
rect 295 41 296 42
rect 296 41 297 42
rect 297 41 298 42
rect 298 41 299 42
rect 299 41 300 42
rect 300 41 301 42
rect 301 41 302 42
rect 302 41 303 42
rect 303 41 304 42
rect 304 41 305 42
rect 305 41 306 42
rect 306 41 307 42
rect 307 41 308 42
rect 308 41 309 42
rect 309 41 310 42
rect 310 41 311 42
rect 311 41 312 42
rect 312 41 313 42
rect 313 41 314 42
rect 314 41 315 42
rect 315 41 316 42
rect 316 41 317 42
rect 317 41 318 42
rect 318 41 319 42
rect 319 41 320 42
rect 320 41 321 42
rect 321 41 322 42
rect 322 41 323 42
rect 323 41 324 42
rect 366 41 367 42
rect 367 41 368 42
rect 368 41 369 42
rect 369 41 370 42
rect 370 41 371 42
rect 371 41 372 42
rect 372 41 373 42
rect 373 41 374 42
rect 374 41 375 42
rect 375 41 376 42
rect 376 41 377 42
rect 377 41 378 42
rect 378 41 379 42
rect 379 41 380 42
rect 214 40 215 41
rect 215 40 216 41
rect 216 40 217 41
rect 255 40 256 41
rect 256 40 257 41
rect 257 40 258 41
rect 258 40 259 41
rect 259 40 260 41
rect 260 40 261 41
rect 261 40 262 41
rect 262 40 263 41
rect 263 40 264 41
rect 264 40 265 41
rect 265 40 266 41
rect 266 40 267 41
rect 267 40 268 41
rect 268 40 269 41
rect 269 40 270 41
rect 270 40 271 41
rect 271 40 272 41
rect 272 40 273 41
rect 273 40 274 41
rect 274 40 275 41
rect 275 40 276 41
rect 276 40 277 41
rect 277 40 278 41
rect 278 40 279 41
rect 279 40 280 41
rect 280 40 281 41
rect 281 40 282 41
rect 282 40 283 41
rect 283 40 284 41
rect 284 40 285 41
rect 285 40 286 41
rect 286 40 287 41
rect 287 40 288 41
rect 288 40 289 41
rect 289 40 290 41
rect 290 40 291 41
rect 291 40 292 41
rect 292 40 293 41
rect 293 40 294 41
rect 294 40 295 41
rect 295 40 296 41
rect 296 40 297 41
rect 297 40 298 41
rect 298 40 299 41
rect 299 40 300 41
rect 300 40 301 41
rect 301 40 302 41
rect 302 40 303 41
rect 303 40 304 41
rect 304 40 305 41
rect 305 40 306 41
rect 306 40 307 41
rect 307 40 308 41
rect 308 40 309 41
rect 309 40 310 41
rect 310 40 311 41
rect 311 40 312 41
rect 312 40 313 41
rect 313 40 314 41
rect 314 40 315 41
rect 315 40 316 41
rect 316 40 317 41
rect 317 40 318 41
rect 318 40 319 41
rect 319 40 320 41
rect 320 40 321 41
rect 321 40 322 41
rect 322 40 323 41
rect 323 40 324 41
rect 324 40 325 41
rect 325 40 326 41
rect 326 40 327 41
rect 327 40 328 41
rect 328 40 329 41
rect 358 40 359 41
rect 359 40 360 41
rect 360 40 361 41
rect 361 40 362 41
rect 362 40 363 41
rect 363 40 364 41
rect 364 40 365 41
rect 365 40 366 41
rect 366 40 367 41
rect 367 40 368 41
rect 368 40 369 41
rect 369 40 370 41
rect 370 40 371 41
rect 371 40 372 41
rect 372 40 373 41
rect 373 40 374 41
rect 374 40 375 41
rect 375 40 376 41
rect 376 40 377 41
rect 377 40 378 41
rect 378 40 379 41
rect 379 40 380 41
rect 263 39 264 40
rect 264 39 265 40
rect 265 39 266 40
rect 266 39 267 40
rect 267 39 268 40
rect 268 39 269 40
rect 269 39 270 40
rect 270 39 271 40
rect 271 39 272 40
rect 272 39 273 40
rect 273 39 274 40
rect 274 39 275 40
rect 275 39 276 40
rect 276 39 277 40
rect 277 39 278 40
rect 278 39 279 40
rect 279 39 280 40
rect 280 39 281 40
rect 281 39 282 40
rect 282 39 283 40
rect 283 39 284 40
rect 284 39 285 40
rect 285 39 286 40
rect 286 39 287 40
rect 287 39 288 40
rect 288 39 289 40
rect 289 39 290 40
rect 290 39 291 40
rect 291 39 292 40
rect 292 39 293 40
rect 293 39 294 40
rect 294 39 295 40
rect 295 39 296 40
rect 296 39 297 40
rect 297 39 298 40
rect 298 39 299 40
rect 299 39 300 40
rect 300 39 301 40
rect 301 39 302 40
rect 302 39 303 40
rect 303 39 304 40
rect 304 39 305 40
rect 305 39 306 40
rect 306 39 307 40
rect 307 39 308 40
rect 308 39 309 40
rect 309 39 310 40
rect 310 39 311 40
rect 311 39 312 40
rect 312 39 313 40
rect 313 39 314 40
rect 314 39 315 40
rect 315 39 316 40
rect 316 39 317 40
rect 317 39 318 40
rect 318 39 319 40
rect 319 39 320 40
rect 320 39 321 40
rect 321 39 322 40
rect 322 39 323 40
rect 323 39 324 40
rect 324 39 325 40
rect 325 39 326 40
rect 326 39 327 40
rect 327 39 328 40
rect 328 39 329 40
rect 358 39 359 40
rect 359 39 360 40
rect 360 39 361 40
rect 361 39 362 40
rect 362 39 363 40
rect 363 39 364 40
rect 364 39 365 40
rect 365 39 366 40
rect 366 39 367 40
rect 367 39 368 40
rect 368 39 369 40
rect 369 39 370 40
rect 370 39 371 40
rect 371 39 372 40
rect 372 39 373 40
rect 373 39 374 40
rect 374 39 375 40
rect 375 39 376 40
rect 376 39 377 40
rect 377 39 378 40
rect 263 38 264 39
rect 264 38 265 39
rect 265 38 266 39
rect 266 38 267 39
rect 267 38 268 39
rect 268 38 269 39
rect 269 38 270 39
rect 270 38 271 39
rect 271 38 272 39
rect 272 38 273 39
rect 273 38 274 39
rect 274 38 275 39
rect 275 38 276 39
rect 276 38 277 39
rect 277 38 278 39
rect 278 38 279 39
rect 279 38 280 39
rect 280 38 281 39
rect 281 38 282 39
rect 282 38 283 39
rect 283 38 284 39
rect 284 38 285 39
rect 285 38 286 39
rect 286 38 287 39
rect 287 38 288 39
rect 288 38 289 39
rect 289 38 290 39
rect 290 38 291 39
rect 291 38 292 39
rect 292 38 293 39
rect 293 38 294 39
rect 294 38 295 39
rect 295 38 296 39
rect 296 38 297 39
rect 297 38 298 39
rect 298 38 299 39
rect 299 38 300 39
rect 300 38 301 39
rect 301 38 302 39
rect 302 38 303 39
rect 303 38 304 39
rect 304 38 305 39
rect 305 38 306 39
rect 306 38 307 39
rect 307 38 308 39
rect 308 38 309 39
rect 309 38 310 39
rect 310 38 311 39
rect 311 38 312 39
rect 312 38 313 39
rect 313 38 314 39
rect 314 38 315 39
rect 315 38 316 39
rect 316 38 317 39
rect 317 38 318 39
rect 318 38 319 39
rect 319 38 320 39
rect 320 38 321 39
rect 321 38 322 39
rect 322 38 323 39
rect 323 38 324 39
rect 324 38 325 39
rect 325 38 326 39
rect 326 38 327 39
rect 327 38 328 39
rect 328 38 329 39
rect 329 38 330 39
rect 330 38 331 39
rect 331 38 332 39
rect 332 38 333 39
rect 333 38 334 39
rect 334 38 335 39
rect 335 38 336 39
rect 336 38 337 39
rect 338 38 339 39
rect 339 38 340 39
rect 340 38 341 39
rect 341 38 342 39
rect 349 38 350 39
rect 350 38 351 39
rect 351 38 352 39
rect 352 38 353 39
rect 353 38 354 39
rect 354 38 355 39
rect 355 38 356 39
rect 356 38 357 39
rect 357 38 358 39
rect 358 38 359 39
rect 359 38 360 39
rect 360 38 361 39
rect 361 38 362 39
rect 362 38 363 39
rect 363 38 364 39
rect 364 38 365 39
rect 365 38 366 39
rect 366 38 367 39
rect 367 38 368 39
rect 368 38 369 39
rect 369 38 370 39
rect 370 38 371 39
rect 371 38 372 39
rect 372 38 373 39
rect 373 38 374 39
rect 374 38 375 39
rect 375 38 376 39
rect 376 38 377 39
rect 377 38 378 39
rect 270 37 271 38
rect 271 37 272 38
rect 272 37 273 38
rect 273 37 274 38
rect 274 37 275 38
rect 275 37 276 38
rect 276 37 277 38
rect 277 37 278 38
rect 278 37 279 38
rect 279 37 280 38
rect 280 37 281 38
rect 281 37 282 38
rect 282 37 283 38
rect 283 37 284 38
rect 284 37 285 38
rect 285 37 286 38
rect 286 37 287 38
rect 287 37 288 38
rect 288 37 289 38
rect 289 37 290 38
rect 290 37 291 38
rect 291 37 292 38
rect 292 37 293 38
rect 293 37 294 38
rect 294 37 295 38
rect 295 37 296 38
rect 296 37 297 38
rect 297 37 298 38
rect 298 37 299 38
rect 299 37 300 38
rect 300 37 301 38
rect 301 37 302 38
rect 302 37 303 38
rect 303 37 304 38
rect 304 37 305 38
rect 305 37 306 38
rect 306 37 307 38
rect 307 37 308 38
rect 308 37 309 38
rect 309 37 310 38
rect 310 37 311 38
rect 311 37 312 38
rect 312 37 313 38
rect 313 37 314 38
rect 314 37 315 38
rect 315 37 316 38
rect 316 37 317 38
rect 317 37 318 38
rect 318 37 319 38
rect 319 37 320 38
rect 320 37 321 38
rect 321 37 322 38
rect 322 37 323 38
rect 323 37 324 38
rect 324 37 325 38
rect 325 37 326 38
rect 326 37 327 38
rect 327 37 328 38
rect 328 37 329 38
rect 329 37 330 38
rect 330 37 331 38
rect 331 37 332 38
rect 332 37 333 38
rect 333 37 334 38
rect 334 37 335 38
rect 335 37 336 38
rect 336 37 337 38
rect 338 37 339 38
rect 339 37 340 38
rect 340 37 341 38
rect 341 37 342 38
rect 349 37 350 38
rect 350 37 351 38
rect 351 37 352 38
rect 352 37 353 38
rect 353 37 354 38
rect 354 37 355 38
rect 355 37 356 38
rect 356 37 357 38
rect 357 37 358 38
rect 358 37 359 38
rect 359 37 360 38
rect 360 37 361 38
rect 361 37 362 38
rect 362 37 363 38
rect 363 37 364 38
rect 364 37 365 38
rect 365 37 366 38
rect 366 37 367 38
rect 367 37 368 38
rect 368 37 369 38
rect 369 37 370 38
rect 370 37 371 38
rect 371 37 372 38
rect 372 37 373 38
rect 373 37 374 38
rect 374 37 375 38
rect 375 37 376 38
rect 270 36 271 37
rect 271 36 272 37
rect 272 36 273 37
rect 273 36 274 37
rect 274 36 275 37
rect 275 36 276 37
rect 276 36 277 37
rect 277 36 278 37
rect 278 36 279 37
rect 279 36 280 37
rect 280 36 281 37
rect 281 36 282 37
rect 282 36 283 37
rect 283 36 284 37
rect 284 36 285 37
rect 285 36 286 37
rect 286 36 287 37
rect 287 36 288 37
rect 288 36 289 37
rect 289 36 290 37
rect 290 36 291 37
rect 291 36 292 37
rect 292 36 293 37
rect 293 36 294 37
rect 294 36 295 37
rect 295 36 296 37
rect 296 36 297 37
rect 297 36 298 37
rect 298 36 299 37
rect 299 36 300 37
rect 300 36 301 37
rect 301 36 302 37
rect 302 36 303 37
rect 303 36 304 37
rect 304 36 305 37
rect 305 36 306 37
rect 306 36 307 37
rect 307 36 308 37
rect 308 36 309 37
rect 309 36 310 37
rect 310 36 311 37
rect 311 36 312 37
rect 312 36 313 37
rect 313 36 314 37
rect 314 36 315 37
rect 315 36 316 37
rect 316 36 317 37
rect 317 36 318 37
rect 318 36 319 37
rect 319 36 320 37
rect 320 36 321 37
rect 321 36 322 37
rect 322 36 323 37
rect 323 36 324 37
rect 324 36 325 37
rect 325 36 326 37
rect 326 36 327 37
rect 327 36 328 37
rect 328 36 329 37
rect 329 36 330 37
rect 330 36 331 37
rect 331 36 332 37
rect 332 36 333 37
rect 333 36 334 37
rect 334 36 335 37
rect 335 36 336 37
rect 336 36 337 37
rect 337 36 338 37
rect 338 36 339 37
rect 339 36 340 37
rect 340 36 341 37
rect 341 36 342 37
rect 342 36 343 37
rect 343 36 344 37
rect 344 36 345 37
rect 345 36 346 37
rect 346 36 347 37
rect 347 36 348 37
rect 348 36 349 37
rect 349 36 350 37
rect 350 36 351 37
rect 351 36 352 37
rect 352 36 353 37
rect 353 36 354 37
rect 354 36 355 37
rect 355 36 356 37
rect 356 36 357 37
rect 357 36 358 37
rect 358 36 359 37
rect 359 36 360 37
rect 360 36 361 37
rect 361 36 362 37
rect 362 36 363 37
rect 363 36 364 37
rect 364 36 365 37
rect 365 36 366 37
rect 366 36 367 37
rect 367 36 368 37
rect 368 36 369 37
rect 369 36 370 37
rect 370 36 371 37
rect 371 36 372 37
rect 372 36 373 37
rect 373 36 374 37
rect 374 36 375 37
rect 375 36 376 37
rect 276 35 277 36
rect 277 35 278 36
rect 278 35 279 36
rect 279 35 280 36
rect 280 35 281 36
rect 281 35 282 36
rect 282 35 283 36
rect 283 35 284 36
rect 284 35 285 36
rect 285 35 286 36
rect 286 35 287 36
rect 287 35 288 36
rect 288 35 289 36
rect 289 35 290 36
rect 290 35 291 36
rect 291 35 292 36
rect 292 35 293 36
rect 293 35 294 36
rect 294 35 295 36
rect 295 35 296 36
rect 296 35 297 36
rect 297 35 298 36
rect 298 35 299 36
rect 299 35 300 36
rect 300 35 301 36
rect 301 35 302 36
rect 302 35 303 36
rect 303 35 304 36
rect 304 35 305 36
rect 305 35 306 36
rect 306 35 307 36
rect 307 35 308 36
rect 308 35 309 36
rect 309 35 310 36
rect 310 35 311 36
rect 311 35 312 36
rect 312 35 313 36
rect 313 35 314 36
rect 314 35 315 36
rect 315 35 316 36
rect 316 35 317 36
rect 317 35 318 36
rect 318 35 319 36
rect 319 35 320 36
rect 320 35 321 36
rect 321 35 322 36
rect 322 35 323 36
rect 323 35 324 36
rect 324 35 325 36
rect 325 35 326 36
rect 326 35 327 36
rect 327 35 328 36
rect 328 35 329 36
rect 329 35 330 36
rect 330 35 331 36
rect 331 35 332 36
rect 332 35 333 36
rect 333 35 334 36
rect 334 35 335 36
rect 335 35 336 36
rect 336 35 337 36
rect 337 35 338 36
rect 338 35 339 36
rect 339 35 340 36
rect 340 35 341 36
rect 341 35 342 36
rect 342 35 343 36
rect 343 35 344 36
rect 344 35 345 36
rect 345 35 346 36
rect 346 35 347 36
rect 347 35 348 36
rect 348 35 349 36
rect 349 35 350 36
rect 350 35 351 36
rect 351 35 352 36
rect 352 35 353 36
rect 353 35 354 36
rect 354 35 355 36
rect 355 35 356 36
rect 356 35 357 36
rect 357 35 358 36
rect 358 35 359 36
rect 359 35 360 36
rect 360 35 361 36
rect 361 35 362 36
rect 362 35 363 36
rect 363 35 364 36
rect 364 35 365 36
rect 365 35 366 36
rect 366 35 367 36
rect 367 35 368 36
rect 368 35 369 36
rect 369 35 370 36
rect 370 35 371 36
rect 371 35 372 36
rect 276 34 277 35
rect 277 34 278 35
rect 278 34 279 35
rect 279 34 280 35
rect 280 34 281 35
rect 281 34 282 35
rect 282 34 283 35
rect 283 34 284 35
rect 284 34 285 35
rect 285 34 286 35
rect 286 34 287 35
rect 287 34 288 35
rect 288 34 289 35
rect 289 34 290 35
rect 290 34 291 35
rect 291 34 292 35
rect 292 34 293 35
rect 293 34 294 35
rect 294 34 295 35
rect 295 34 296 35
rect 296 34 297 35
rect 297 34 298 35
rect 298 34 299 35
rect 299 34 300 35
rect 300 34 301 35
rect 301 34 302 35
rect 302 34 303 35
rect 303 34 304 35
rect 304 34 305 35
rect 305 34 306 35
rect 306 34 307 35
rect 307 34 308 35
rect 308 34 309 35
rect 309 34 310 35
rect 310 34 311 35
rect 311 34 312 35
rect 312 34 313 35
rect 313 34 314 35
rect 314 34 315 35
rect 315 34 316 35
rect 316 34 317 35
rect 317 34 318 35
rect 318 34 319 35
rect 319 34 320 35
rect 320 34 321 35
rect 321 34 322 35
rect 322 34 323 35
rect 323 34 324 35
rect 324 34 325 35
rect 325 34 326 35
rect 326 34 327 35
rect 327 34 328 35
rect 328 34 329 35
rect 329 34 330 35
rect 330 34 331 35
rect 331 34 332 35
rect 332 34 333 35
rect 333 34 334 35
rect 334 34 335 35
rect 335 34 336 35
rect 336 34 337 35
rect 337 34 338 35
rect 338 34 339 35
rect 339 34 340 35
rect 340 34 341 35
rect 341 34 342 35
rect 342 34 343 35
rect 343 34 344 35
rect 344 34 345 35
rect 345 34 346 35
rect 346 34 347 35
rect 347 34 348 35
rect 348 34 349 35
rect 349 34 350 35
rect 350 34 351 35
rect 351 34 352 35
rect 352 34 353 35
rect 353 34 354 35
rect 354 34 355 35
rect 355 34 356 35
rect 356 34 357 35
rect 357 34 358 35
rect 358 34 359 35
rect 359 34 360 35
rect 360 34 361 35
rect 361 34 362 35
rect 362 34 363 35
rect 363 34 364 35
rect 364 34 365 35
rect 365 34 366 35
rect 366 34 367 35
rect 367 34 368 35
rect 368 34 369 35
rect 369 34 370 35
rect 370 34 371 35
rect 371 34 372 35
rect 281 33 282 34
rect 282 33 283 34
rect 283 33 284 34
rect 284 33 285 34
rect 285 33 286 34
rect 286 33 287 34
rect 287 33 288 34
rect 288 33 289 34
rect 289 33 290 34
rect 290 33 291 34
rect 291 33 292 34
rect 292 33 293 34
rect 293 33 294 34
rect 294 33 295 34
rect 295 33 296 34
rect 296 33 297 34
rect 297 33 298 34
rect 298 33 299 34
rect 299 33 300 34
rect 300 33 301 34
rect 301 33 302 34
rect 302 33 303 34
rect 303 33 304 34
rect 304 33 305 34
rect 305 33 306 34
rect 306 33 307 34
rect 307 33 308 34
rect 308 33 309 34
rect 309 33 310 34
rect 310 33 311 34
rect 311 33 312 34
rect 312 33 313 34
rect 313 33 314 34
rect 314 33 315 34
rect 315 33 316 34
rect 316 33 317 34
rect 317 33 318 34
rect 318 33 319 34
rect 319 33 320 34
rect 320 33 321 34
rect 321 33 322 34
rect 322 33 323 34
rect 323 33 324 34
rect 324 33 325 34
rect 325 33 326 34
rect 326 33 327 34
rect 327 33 328 34
rect 328 33 329 34
rect 329 33 330 34
rect 330 33 331 34
rect 331 33 332 34
rect 332 33 333 34
rect 333 33 334 34
rect 334 33 335 34
rect 335 33 336 34
rect 336 33 337 34
rect 337 33 338 34
rect 338 33 339 34
rect 339 33 340 34
rect 340 33 341 34
rect 341 33 342 34
rect 342 33 343 34
rect 343 33 344 34
rect 344 33 345 34
rect 345 33 346 34
rect 346 33 347 34
rect 347 33 348 34
rect 348 33 349 34
rect 349 33 350 34
rect 350 33 351 34
rect 351 33 352 34
rect 352 33 353 34
rect 353 33 354 34
rect 354 33 355 34
rect 355 33 356 34
rect 356 33 357 34
rect 357 33 358 34
rect 358 33 359 34
rect 359 33 360 34
rect 360 33 361 34
rect 361 33 362 34
rect 362 33 363 34
rect 363 33 364 34
rect 364 33 365 34
rect 365 33 366 34
rect 366 33 367 34
rect 367 33 368 34
rect 368 33 369 34
rect 369 33 370 34
rect 281 32 282 33
rect 282 32 283 33
rect 283 32 284 33
rect 284 32 285 33
rect 285 32 286 33
rect 286 32 287 33
rect 287 32 288 33
rect 288 32 289 33
rect 289 32 290 33
rect 290 32 291 33
rect 291 32 292 33
rect 292 32 293 33
rect 293 32 294 33
rect 294 32 295 33
rect 295 32 296 33
rect 296 32 297 33
rect 297 32 298 33
rect 298 32 299 33
rect 299 32 300 33
rect 300 32 301 33
rect 301 32 302 33
rect 302 32 303 33
rect 303 32 304 33
rect 304 32 305 33
rect 305 32 306 33
rect 306 32 307 33
rect 307 32 308 33
rect 308 32 309 33
rect 309 32 310 33
rect 310 32 311 33
rect 311 32 312 33
rect 312 32 313 33
rect 313 32 314 33
rect 314 32 315 33
rect 315 32 316 33
rect 316 32 317 33
rect 317 32 318 33
rect 318 32 319 33
rect 319 32 320 33
rect 320 32 321 33
rect 321 32 322 33
rect 322 32 323 33
rect 323 32 324 33
rect 324 32 325 33
rect 325 32 326 33
rect 326 32 327 33
rect 327 32 328 33
rect 328 32 329 33
rect 329 32 330 33
rect 330 32 331 33
rect 331 32 332 33
rect 332 32 333 33
rect 333 32 334 33
rect 334 32 335 33
rect 335 32 336 33
rect 336 32 337 33
rect 337 32 338 33
rect 338 32 339 33
rect 339 32 340 33
rect 340 32 341 33
rect 341 32 342 33
rect 342 32 343 33
rect 343 32 344 33
rect 344 32 345 33
rect 345 32 346 33
rect 346 32 347 33
rect 347 32 348 33
rect 348 32 349 33
rect 349 32 350 33
rect 350 32 351 33
rect 351 32 352 33
rect 352 32 353 33
rect 353 32 354 33
rect 354 32 355 33
rect 355 32 356 33
rect 356 32 357 33
rect 357 32 358 33
rect 358 32 359 33
rect 359 32 360 33
rect 360 32 361 33
rect 361 32 362 33
rect 362 32 363 33
rect 363 32 364 33
rect 364 32 365 33
rect 365 32 366 33
rect 366 32 367 33
rect 367 32 368 33
rect 368 32 369 33
rect 369 32 370 33
rect 287 31 288 32
rect 288 31 289 32
rect 289 31 290 32
rect 290 31 291 32
rect 291 31 292 32
rect 292 31 293 32
rect 293 31 294 32
rect 294 31 295 32
rect 295 31 296 32
rect 296 31 297 32
rect 297 31 298 32
rect 298 31 299 32
rect 299 31 300 32
rect 300 31 301 32
rect 301 31 302 32
rect 302 31 303 32
rect 303 31 304 32
rect 304 31 305 32
rect 305 31 306 32
rect 306 31 307 32
rect 307 31 308 32
rect 308 31 309 32
rect 309 31 310 32
rect 310 31 311 32
rect 311 31 312 32
rect 312 31 313 32
rect 313 31 314 32
rect 314 31 315 32
rect 315 31 316 32
rect 316 31 317 32
rect 317 31 318 32
rect 318 31 319 32
rect 319 31 320 32
rect 320 31 321 32
rect 321 31 322 32
rect 322 31 323 32
rect 323 31 324 32
rect 324 31 325 32
rect 325 31 326 32
rect 326 31 327 32
rect 327 31 328 32
rect 328 31 329 32
rect 329 31 330 32
rect 330 31 331 32
rect 331 31 332 32
rect 332 31 333 32
rect 333 31 334 32
rect 334 31 335 32
rect 335 31 336 32
rect 336 31 337 32
rect 337 31 338 32
rect 338 31 339 32
rect 339 31 340 32
rect 340 31 341 32
rect 341 31 342 32
rect 342 31 343 32
rect 343 31 344 32
rect 344 31 345 32
rect 345 31 346 32
rect 346 31 347 32
rect 347 31 348 32
rect 348 31 349 32
rect 349 31 350 32
rect 350 31 351 32
rect 351 31 352 32
rect 352 31 353 32
rect 353 31 354 32
rect 354 31 355 32
rect 355 31 356 32
rect 356 31 357 32
rect 357 31 358 32
rect 358 31 359 32
rect 359 31 360 32
rect 360 31 361 32
rect 361 31 362 32
rect 362 31 363 32
rect 363 31 364 32
rect 364 31 365 32
rect 365 31 366 32
rect 366 31 367 32
rect 287 30 288 31
rect 288 30 289 31
rect 289 30 290 31
rect 290 30 291 31
rect 291 30 292 31
rect 292 30 293 31
rect 293 30 294 31
rect 294 30 295 31
rect 295 30 296 31
rect 296 30 297 31
rect 297 30 298 31
rect 298 30 299 31
rect 299 30 300 31
rect 300 30 301 31
rect 301 30 302 31
rect 302 30 303 31
rect 303 30 304 31
rect 304 30 305 31
rect 305 30 306 31
rect 306 30 307 31
rect 307 30 308 31
rect 308 30 309 31
rect 309 30 310 31
rect 310 30 311 31
rect 311 30 312 31
rect 312 30 313 31
rect 313 30 314 31
rect 314 30 315 31
rect 315 30 316 31
rect 316 30 317 31
rect 317 30 318 31
rect 318 30 319 31
rect 319 30 320 31
rect 320 30 321 31
rect 321 30 322 31
rect 322 30 323 31
rect 323 30 324 31
rect 324 30 325 31
rect 325 30 326 31
rect 326 30 327 31
rect 327 30 328 31
rect 328 30 329 31
rect 329 30 330 31
rect 330 30 331 31
rect 331 30 332 31
rect 332 30 333 31
rect 333 30 334 31
rect 334 30 335 31
rect 335 30 336 31
rect 336 30 337 31
rect 337 30 338 31
rect 338 30 339 31
rect 339 30 340 31
rect 340 30 341 31
rect 341 30 342 31
rect 342 30 343 31
rect 343 30 344 31
rect 344 30 345 31
rect 345 30 346 31
rect 346 30 347 31
rect 347 30 348 31
rect 348 30 349 31
rect 349 30 350 31
rect 350 30 351 31
rect 351 30 352 31
rect 352 30 353 31
rect 353 30 354 31
rect 354 30 355 31
rect 355 30 356 31
rect 356 30 357 31
rect 357 30 358 31
rect 358 30 359 31
rect 359 30 360 31
rect 360 30 361 31
rect 361 30 362 31
rect 362 30 363 31
rect 363 30 364 31
rect 364 30 365 31
rect 365 30 366 31
rect 366 30 367 31
rect 293 29 294 30
rect 294 29 295 30
rect 295 29 296 30
rect 296 29 297 30
rect 297 29 298 30
rect 298 29 299 30
rect 299 29 300 30
rect 300 29 301 30
rect 301 29 302 30
rect 302 29 303 30
rect 303 29 304 30
rect 304 29 305 30
rect 305 29 306 30
rect 306 29 307 30
rect 307 29 308 30
rect 308 29 309 30
rect 309 29 310 30
rect 310 29 311 30
rect 311 29 312 30
rect 312 29 313 30
rect 313 29 314 30
rect 314 29 315 30
rect 315 29 316 30
rect 316 29 317 30
rect 317 29 318 30
rect 318 29 319 30
rect 319 29 320 30
rect 320 29 321 30
rect 321 29 322 30
rect 322 29 323 30
rect 323 29 324 30
rect 324 29 325 30
rect 325 29 326 30
rect 326 29 327 30
rect 327 29 328 30
rect 328 29 329 30
rect 329 29 330 30
rect 330 29 331 30
rect 331 29 332 30
rect 332 29 333 30
rect 333 29 334 30
rect 334 29 335 30
rect 335 29 336 30
rect 336 29 337 30
rect 337 29 338 30
rect 338 29 339 30
rect 339 29 340 30
rect 340 29 341 30
rect 341 29 342 30
rect 342 29 343 30
rect 343 29 344 30
rect 344 29 345 30
rect 345 29 346 30
rect 346 29 347 30
rect 347 29 348 30
rect 348 29 349 30
rect 349 29 350 30
rect 350 29 351 30
rect 351 29 352 30
rect 352 29 353 30
rect 353 29 354 30
rect 354 29 355 30
rect 355 29 356 30
rect 356 29 357 30
rect 357 29 358 30
rect 358 29 359 30
rect 359 29 360 30
rect 360 29 361 30
rect 361 29 362 30
rect 362 29 363 30
rect 363 29 364 30
rect 364 29 365 30
rect 293 28 294 29
rect 294 28 295 29
rect 295 28 296 29
rect 296 28 297 29
rect 297 28 298 29
rect 298 28 299 29
rect 299 28 300 29
rect 300 28 301 29
rect 301 28 302 29
rect 302 28 303 29
rect 303 28 304 29
rect 304 28 305 29
rect 305 28 306 29
rect 306 28 307 29
rect 307 28 308 29
rect 308 28 309 29
rect 309 28 310 29
rect 310 28 311 29
rect 311 28 312 29
rect 312 28 313 29
rect 313 28 314 29
rect 314 28 315 29
rect 315 28 316 29
rect 316 28 317 29
rect 317 28 318 29
rect 318 28 319 29
rect 319 28 320 29
rect 320 28 321 29
rect 321 28 322 29
rect 322 28 323 29
rect 323 28 324 29
rect 324 28 325 29
rect 325 28 326 29
rect 326 28 327 29
rect 327 28 328 29
rect 328 28 329 29
rect 329 28 330 29
rect 330 28 331 29
rect 331 28 332 29
rect 332 28 333 29
rect 333 28 334 29
rect 334 28 335 29
rect 335 28 336 29
rect 336 28 337 29
rect 337 28 338 29
rect 338 28 339 29
rect 339 28 340 29
rect 340 28 341 29
rect 341 28 342 29
rect 342 28 343 29
rect 343 28 344 29
rect 344 28 345 29
rect 345 28 346 29
rect 346 28 347 29
rect 347 28 348 29
rect 348 28 349 29
rect 349 28 350 29
rect 350 28 351 29
rect 351 28 352 29
rect 352 28 353 29
rect 353 28 354 29
rect 354 28 355 29
rect 355 28 356 29
rect 356 28 357 29
rect 357 28 358 29
rect 358 28 359 29
rect 359 28 360 29
rect 360 28 361 29
rect 361 28 362 29
rect 362 28 363 29
rect 363 28 364 29
rect 364 28 365 29
rect 298 27 299 28
rect 299 27 300 28
rect 300 27 301 28
rect 301 27 302 28
rect 302 27 303 28
rect 303 27 304 28
rect 304 27 305 28
rect 305 27 306 28
rect 306 27 307 28
rect 307 27 308 28
rect 308 27 309 28
rect 309 27 310 28
rect 310 27 311 28
rect 311 27 312 28
rect 312 27 313 28
rect 313 27 314 28
rect 314 27 315 28
rect 315 27 316 28
rect 316 27 317 28
rect 317 27 318 28
rect 318 27 319 28
rect 319 27 320 28
rect 320 27 321 28
rect 321 27 322 28
rect 322 27 323 28
rect 323 27 324 28
rect 324 27 325 28
rect 325 27 326 28
rect 326 27 327 28
rect 327 27 328 28
rect 328 27 329 28
rect 329 27 330 28
rect 330 27 331 28
rect 331 27 332 28
rect 332 27 333 28
rect 333 27 334 28
rect 334 27 335 28
rect 335 27 336 28
rect 336 27 337 28
rect 337 27 338 28
rect 338 27 339 28
rect 339 27 340 28
rect 340 27 341 28
rect 341 27 342 28
rect 342 27 343 28
rect 343 27 344 28
rect 344 27 345 28
rect 345 27 346 28
rect 346 27 347 28
rect 347 27 348 28
rect 348 27 349 28
rect 349 27 350 28
rect 350 27 351 28
rect 351 27 352 28
rect 352 27 353 28
rect 353 27 354 28
rect 354 27 355 28
rect 355 27 356 28
rect 356 27 357 28
rect 357 27 358 28
rect 358 27 359 28
rect 359 27 360 28
rect 360 27 361 28
rect 298 26 299 27
rect 299 26 300 27
rect 300 26 301 27
rect 301 26 302 27
rect 302 26 303 27
rect 303 26 304 27
rect 304 26 305 27
rect 305 26 306 27
rect 306 26 307 27
rect 307 26 308 27
rect 308 26 309 27
rect 309 26 310 27
rect 310 26 311 27
rect 311 26 312 27
rect 312 26 313 27
rect 313 26 314 27
rect 314 26 315 27
rect 315 26 316 27
rect 316 26 317 27
rect 317 26 318 27
rect 318 26 319 27
rect 319 26 320 27
rect 320 26 321 27
rect 321 26 322 27
rect 322 26 323 27
rect 323 26 324 27
rect 324 26 325 27
rect 325 26 326 27
rect 326 26 327 27
rect 327 26 328 27
rect 328 26 329 27
rect 329 26 330 27
rect 330 26 331 27
rect 331 26 332 27
rect 332 26 333 27
rect 333 26 334 27
rect 334 26 335 27
rect 335 26 336 27
rect 336 26 337 27
rect 337 26 338 27
rect 338 26 339 27
rect 339 26 340 27
rect 340 26 341 27
rect 341 26 342 27
rect 342 26 343 27
rect 343 26 344 27
rect 344 26 345 27
rect 345 26 346 27
rect 346 26 347 27
rect 347 26 348 27
rect 348 26 349 27
rect 349 26 350 27
rect 350 26 351 27
rect 351 26 352 27
rect 352 26 353 27
rect 353 26 354 27
rect 354 26 355 27
rect 355 26 356 27
rect 356 26 357 27
rect 357 26 358 27
rect 358 26 359 27
rect 359 26 360 27
rect 360 26 361 27
rect 298 25 299 26
rect 299 25 300 26
rect 300 25 301 26
rect 301 25 302 26
rect 302 25 303 26
rect 303 25 304 26
rect 304 25 305 26
rect 305 25 306 26
rect 306 25 307 26
rect 307 25 308 26
rect 308 25 309 26
rect 309 25 310 26
rect 310 25 311 26
rect 311 25 312 26
rect 312 25 313 26
rect 313 25 314 26
rect 314 25 315 26
rect 315 25 316 26
rect 316 25 317 26
rect 317 25 318 26
rect 318 25 319 26
rect 319 25 320 26
rect 320 25 321 26
rect 321 25 322 26
rect 322 25 323 26
rect 323 25 324 26
rect 324 25 325 26
rect 325 25 326 26
rect 326 25 327 26
rect 327 25 328 26
rect 328 25 329 26
rect 329 25 330 26
rect 330 25 331 26
rect 331 25 332 26
rect 332 25 333 26
rect 333 25 334 26
rect 334 25 335 26
rect 335 25 336 26
rect 336 25 337 26
rect 337 25 338 26
rect 338 25 339 26
rect 339 25 340 26
rect 340 25 341 26
rect 341 25 342 26
rect 342 25 343 26
rect 343 25 344 26
rect 344 25 345 26
rect 345 25 346 26
rect 346 25 347 26
rect 347 25 348 26
rect 348 25 349 26
rect 349 25 350 26
rect 350 25 351 26
rect 351 25 352 26
rect 352 25 353 26
rect 353 25 354 26
rect 354 25 355 26
rect 355 25 356 26
rect 356 25 357 26
rect 357 25 358 26
rect 358 25 359 26
rect 359 25 360 26
rect 360 25 361 26
rect 304 24 305 25
rect 305 24 306 25
rect 306 24 307 25
rect 307 24 308 25
rect 308 24 309 25
rect 309 24 310 25
rect 310 24 311 25
rect 311 24 312 25
rect 312 24 313 25
rect 313 24 314 25
rect 314 24 315 25
rect 315 24 316 25
rect 316 24 317 25
rect 317 24 318 25
rect 318 24 319 25
rect 319 24 320 25
rect 320 24 321 25
rect 321 24 322 25
rect 322 24 323 25
rect 323 24 324 25
rect 324 24 325 25
rect 325 24 326 25
rect 326 24 327 25
rect 327 24 328 25
rect 328 24 329 25
rect 329 24 330 25
rect 330 24 331 25
rect 331 24 332 25
rect 332 24 333 25
rect 333 24 334 25
rect 334 24 335 25
rect 335 24 336 25
rect 336 24 337 25
rect 337 24 338 25
rect 338 24 339 25
rect 339 24 340 25
rect 340 24 341 25
rect 341 24 342 25
rect 342 24 343 25
rect 343 24 344 25
rect 344 24 345 25
rect 345 24 346 25
rect 346 24 347 25
rect 347 24 348 25
rect 348 24 349 25
rect 349 24 350 25
rect 350 24 351 25
rect 351 24 352 25
rect 352 24 353 25
rect 353 24 354 25
rect 354 24 355 25
rect 355 24 356 25
rect 356 24 357 25
rect 357 24 358 25
rect 358 24 359 25
rect 304 23 305 24
rect 305 23 306 24
rect 306 23 307 24
rect 307 23 308 24
rect 308 23 309 24
rect 309 23 310 24
rect 310 23 311 24
rect 311 23 312 24
rect 312 23 313 24
rect 313 23 314 24
rect 314 23 315 24
rect 315 23 316 24
rect 316 23 317 24
rect 317 23 318 24
rect 318 23 319 24
rect 319 23 320 24
rect 320 23 321 24
rect 321 23 322 24
rect 322 23 323 24
rect 323 23 324 24
rect 324 23 325 24
rect 325 23 326 24
rect 326 23 327 24
rect 327 23 328 24
rect 328 23 329 24
rect 329 23 330 24
rect 330 23 331 24
rect 331 23 332 24
rect 332 23 333 24
rect 333 23 334 24
rect 334 23 335 24
rect 335 23 336 24
rect 336 23 337 24
rect 337 23 338 24
rect 338 23 339 24
rect 339 23 340 24
rect 340 23 341 24
rect 341 23 342 24
rect 342 23 343 24
rect 343 23 344 24
rect 344 23 345 24
rect 345 23 346 24
rect 346 23 347 24
rect 347 23 348 24
rect 348 23 349 24
rect 349 23 350 24
rect 350 23 351 24
rect 351 23 352 24
rect 352 23 353 24
rect 353 23 354 24
rect 354 23 355 24
rect 355 23 356 24
rect 356 23 357 24
rect 357 23 358 24
rect 358 23 359 24
rect 309 22 310 23
rect 310 22 311 23
rect 311 22 312 23
rect 312 22 313 23
rect 313 22 314 23
rect 314 22 315 23
rect 315 22 316 23
rect 316 22 317 23
rect 317 22 318 23
rect 318 22 319 23
rect 319 22 320 23
rect 320 22 321 23
rect 321 22 322 23
rect 322 22 323 23
rect 323 22 324 23
rect 324 22 325 23
rect 325 22 326 23
rect 326 22 327 23
rect 327 22 328 23
rect 328 22 329 23
rect 329 22 330 23
rect 330 22 331 23
rect 331 22 332 23
rect 332 22 333 23
rect 333 22 334 23
rect 334 22 335 23
rect 335 22 336 23
rect 336 22 337 23
rect 337 22 338 23
rect 338 22 339 23
rect 339 22 340 23
rect 340 22 341 23
rect 341 22 342 23
rect 342 22 343 23
rect 343 22 344 23
rect 344 22 345 23
rect 345 22 346 23
rect 346 22 347 23
rect 347 22 348 23
rect 348 22 349 23
rect 349 22 350 23
rect 350 22 351 23
rect 351 22 352 23
rect 352 22 353 23
rect 353 22 354 23
rect 354 22 355 23
rect 355 22 356 23
rect 356 22 357 23
rect 309 21 310 22
rect 310 21 311 22
rect 311 21 312 22
rect 312 21 313 22
rect 313 21 314 22
rect 314 21 315 22
rect 315 21 316 22
rect 316 21 317 22
rect 317 21 318 22
rect 318 21 319 22
rect 319 21 320 22
rect 320 21 321 22
rect 321 21 322 22
rect 322 21 323 22
rect 323 21 324 22
rect 324 21 325 22
rect 325 21 326 22
rect 326 21 327 22
rect 327 21 328 22
rect 328 21 329 22
rect 329 21 330 22
rect 330 21 331 22
rect 331 21 332 22
rect 332 21 333 22
rect 333 21 334 22
rect 334 21 335 22
rect 335 21 336 22
rect 336 21 337 22
rect 337 21 338 22
rect 338 21 339 22
rect 339 21 340 22
rect 340 21 341 22
rect 341 21 342 22
rect 342 21 343 22
rect 343 21 344 22
rect 344 21 345 22
rect 345 21 346 22
rect 346 21 347 22
rect 347 21 348 22
rect 348 21 349 22
rect 349 21 350 22
rect 350 21 351 22
rect 351 21 352 22
rect 352 21 353 22
rect 353 21 354 22
rect 354 21 355 22
rect 355 21 356 22
rect 356 21 357 22
rect 317 20 318 21
rect 318 20 319 21
rect 319 20 320 21
rect 320 20 321 21
rect 321 20 322 21
rect 322 20 323 21
rect 323 20 324 21
rect 324 20 325 21
rect 325 20 326 21
rect 326 20 327 21
rect 327 20 328 21
rect 328 20 329 21
rect 329 20 330 21
rect 330 20 331 21
rect 331 20 332 21
rect 332 20 333 21
rect 333 20 334 21
rect 334 20 335 21
rect 335 20 336 21
rect 336 20 337 21
rect 337 20 338 21
rect 338 20 339 21
rect 339 20 340 21
rect 340 20 341 21
rect 341 20 342 21
rect 342 20 343 21
rect 343 20 344 21
rect 344 20 345 21
rect 345 20 346 21
rect 346 20 347 21
rect 347 20 348 21
rect 348 20 349 21
rect 349 20 350 21
rect 350 20 351 21
rect 351 20 352 21
rect 352 20 353 21
rect 353 20 354 21
rect 317 19 318 20
rect 318 19 319 20
rect 319 19 320 20
rect 320 19 321 20
rect 321 19 322 20
rect 322 19 323 20
rect 323 19 324 20
rect 324 19 325 20
rect 325 19 326 20
rect 326 19 327 20
rect 327 19 328 20
rect 328 19 329 20
rect 329 19 330 20
rect 330 19 331 20
rect 331 19 332 20
rect 332 19 333 20
rect 333 19 334 20
rect 334 19 335 20
rect 335 19 336 20
rect 336 19 337 20
rect 337 19 338 20
rect 338 19 339 20
rect 339 19 340 20
rect 340 19 341 20
rect 341 19 342 20
rect 342 19 343 20
rect 343 19 344 20
rect 344 19 345 20
rect 345 19 346 20
rect 346 19 347 20
rect 347 19 348 20
rect 348 19 349 20
rect 349 19 350 20
rect 350 19 351 20
rect 351 19 352 20
rect 352 19 353 20
rect 353 19 354 20
rect 326 18 327 19
rect 327 18 328 19
rect 328 18 329 19
rect 329 18 330 19
rect 330 18 331 19
rect 331 18 332 19
rect 332 18 333 19
rect 333 18 334 19
rect 334 18 335 19
rect 335 18 336 19
rect 336 18 337 19
rect 337 18 338 19
rect 338 18 339 19
rect 339 18 340 19
rect 340 18 341 19
rect 341 18 342 19
rect 342 18 343 19
rect 343 18 344 19
rect 344 18 345 19
rect 345 18 346 19
rect 346 18 347 19
rect 347 18 348 19
rect 348 18 349 19
rect 349 18 350 19
rect 350 18 351 19
rect 351 18 352 19
rect 326 17 327 18
rect 327 17 328 18
rect 328 17 329 18
rect 329 17 330 18
rect 330 17 331 18
rect 331 17 332 18
rect 332 17 333 18
rect 333 17 334 18
rect 334 17 335 18
rect 335 17 336 18
rect 336 17 337 18
rect 337 17 338 18
rect 338 17 339 18
rect 339 17 340 18
rect 340 17 341 18
rect 341 17 342 18
rect 342 17 343 18
rect 343 17 344 18
rect 344 17 345 18
rect 345 17 346 18
rect 346 17 347 18
rect 347 17 348 18
rect 348 17 349 18
rect 349 17 350 18
rect 350 17 351 18
rect 351 17 352 18
<< end >>
