* Extracted by KLayout

.SUBCKT TOP A Q SUBSTRATE
X$1 \$5 \$1 Q SUBSTRATE INV
X$2 \$5 A \$1 SUBSTRATE INV
.ENDS TOP

.SUBCKT INV \$2 \$4 \$5 SUBSTRATE
M$1 \$2 \$4 \$5 \$2 PMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P PS=3.45U
+ PD=3.45U
M$2 SUBSTRATE \$4 \$5 SUBSTRATE NMOS L=0.25U W=0.95U AS=0.73625P AD=0.73625P
+ PS=3.45U PD=3.45U
.ENDS INV
