magic
tech scmos
timestamp 1537343441
<< metal1 >>
rect 4 96 8 100
rect 92 96 96 100
rect 0 92 100 96
rect 4 84 96 92
rect 4 80 16 84
rect 20 80 24 84
rect 76 80 80 84
rect 84 80 96 84
rect 4 76 96 80
rect 4 24 16 76
rect 20 68 80 76
rect 20 64 32 68
rect 36 64 40 68
rect 60 64 64 68
rect 68 64 80 68
rect 20 60 80 64
rect 20 40 32 60
rect 36 52 64 60
rect 36 48 48 52
rect 52 48 64 52
rect 36 40 64 48
rect 68 40 80 60
rect 20 36 80 40
rect 20 32 32 36
rect 36 32 40 36
rect 60 32 64 36
rect 68 32 80 36
rect 20 24 80 32
rect 84 24 96 76
rect 4 20 96 24
rect 4 16 16 20
rect 20 16 24 20
rect 76 16 80 20
rect 84 16 96 20
rect 4 8 96 16
rect 0 4 100 8
rect 4 0 8 4
rect 92 0 96 4
<< metal2 >>
rect 4 96 8 100
rect 92 96 96 100
rect 0 92 100 96
rect 4 88 8 92
rect 12 88 16 92
rect 84 88 88 92
rect 92 88 96 92
rect 4 84 96 88
rect 4 16 8 84
rect 12 80 16 84
rect 20 80 24 84
rect 76 80 80 84
rect 84 80 88 84
rect 12 76 88 80
rect 12 24 16 76
rect 20 72 24 76
rect 28 72 32 76
rect 68 72 72 76
rect 76 72 80 76
rect 20 68 80 72
rect 20 32 24 68
rect 28 64 32 68
rect 36 64 40 68
rect 60 64 64 68
rect 68 64 72 68
rect 28 60 72 64
rect 28 40 32 60
rect 36 56 40 60
rect 44 56 48 60
rect 52 56 56 60
rect 60 56 64 60
rect 36 52 64 56
rect 36 48 40 52
rect 44 48 48 52
rect 52 48 56 52
rect 60 48 64 52
rect 36 44 64 48
rect 36 40 40 44
rect 44 40 48 44
rect 52 40 56 44
rect 60 40 64 44
rect 68 40 72 60
rect 28 36 72 40
rect 28 32 32 36
rect 36 32 40 36
rect 60 32 64 36
rect 68 32 72 36
rect 76 32 80 68
rect 20 28 80 32
rect 20 24 24 28
rect 28 24 32 28
rect 68 24 72 28
rect 76 24 80 28
rect 84 24 88 76
rect 12 20 88 24
rect 12 16 16 20
rect 20 16 24 20
rect 76 16 80 20
rect 84 16 88 20
rect 92 16 96 84
rect 4 12 96 16
rect 4 8 8 12
rect 12 8 16 12
rect 84 8 88 12
rect 92 8 96 12
rect 0 4 100 8
rect 4 0 8 4
rect 92 0 96 4
<< metal3 >>
rect 0 92 100 100
rect 0 88 8 92
rect 12 88 16 92
rect 84 88 88 92
rect 92 88 100 92
rect 0 84 100 88
rect 0 16 8 84
rect 12 76 88 84
rect 12 72 24 76
rect 28 72 32 76
rect 68 72 72 76
rect 76 72 88 76
rect 12 68 88 72
rect 12 32 24 68
rect 28 60 72 68
rect 28 56 40 60
rect 44 56 48 60
rect 52 56 56 60
rect 60 56 72 60
rect 28 52 72 56
rect 28 48 40 52
rect 44 48 56 52
rect 60 48 72 52
rect 28 44 72 48
rect 28 40 40 44
rect 44 40 48 44
rect 52 40 56 44
rect 60 40 72 44
rect 28 32 72 40
rect 76 32 88 68
rect 12 28 88 32
rect 12 24 24 28
rect 28 24 32 28
rect 68 24 72 28
rect 76 24 88 28
rect 12 16 88 24
rect 92 16 100 84
rect 0 12 100 16
rect 0 8 8 12
rect 12 8 16 12
rect 84 8 88 12
rect 92 8 100 12
rect 0 0 100 8
<< m2contact >>
rect 0 96 4 100
rect 8 96 92 100
rect 96 96 100 100
rect 0 8 4 92
rect 16 80 20 84
rect 24 80 76 84
rect 80 80 84 84
rect 16 24 20 76
rect 32 64 36 68
rect 40 64 60 68
rect 64 64 68 68
rect 32 40 36 60
rect 48 48 52 52
rect 64 40 68 60
rect 32 32 36 36
rect 40 32 60 36
rect 64 32 68 36
rect 80 24 84 76
rect 16 16 20 20
rect 24 16 76 20
rect 80 16 84 20
rect 96 8 100 92
rect 0 0 4 4
rect 8 0 92 4
rect 96 0 100 4
<< m3contact >>
rect 8 88 12 92
rect 16 88 84 92
rect 88 88 92 92
rect 8 16 12 84
rect 24 72 28 76
rect 32 72 68 76
rect 72 72 76 76
rect 24 32 28 68
rect 40 56 44 60
rect 48 56 52 60
rect 56 56 60 60
rect 40 48 44 52
rect 56 48 60 52
rect 40 40 44 44
rect 48 40 52 44
rect 56 40 60 44
rect 72 32 76 68
rect 24 24 28 28
rect 32 24 68 28
rect 72 24 76 28
rect 88 16 92 84
rect 8 8 12 12
rect 16 8 84 12
rect 88 8 92 12
<< glass >>
rect 12 12 88 88
<< end >>
