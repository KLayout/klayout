* Extracted by KLayout

* cell SP6TArray_2X4
.SUBCKT SP6TArray_2X4
* net 1 bl[0]
* net 2 bl_n[0]
* net 3 bl[1]
* net 4 bl_n[1]
* net 5 bl[2]
* net 6 bl_n[2]
* net 7 bl[3]
* net 8 bl_n[3]
* net 9 vdd
* net 10 wl[0]
* net 11 wl[1]
* net 12 vss
* cell instance $1 r0 *1 0,0
X$1 1 2 3 4 9 10 11 12 SP6TArray_2X2
* cell instance $2 r0 *1 4.36,0
X$2 5 6 7 8 9 10 11 12 SP6TArray_2X2
.ENDS SP6TArray_2X4

* cell SP6TArray_2X2
* pin bl[0]
* pin bl_n[0]
* pin bl[1]
* pin bl_n[1]
* pin vdd
* pin wl[0]
* pin wl[1]
* pin vss
.SUBCKT SP6TArray_2X2 1 2 3 4 5 6 7 8
* net 1 bl[0]
* net 2 bl_n[0]
* net 3 bl[1]
* net 4 bl_n[1]
* net 5 vdd
* net 6 wl[0]
* net 7 wl[1]
* net 8 vss
* cell instance $1 r0 *1 0,0
X$1 1 2 5 6 7 8 SP6TArray_2X1
* cell instance $2 r0 *1 2.18,0
X$2 3 4 5 6 7 8 SP6TArray_2X1
.ENDS SP6TArray_2X2

* cell SP6TArray_2X1
* pin bl[0]
* pin bl_n[0]
* pin vdd
* pin wl[0]
* pin wl[1]
* pin vss
.SUBCKT SP6TArray_2X1 1 2 3 4 5 6
* net 1 bl[0]
* net 2 bl_n[0]
* net 3 vdd
* net 4 wl[0]
* net 5 wl[1]
* net 6 vss
* cell instance $1 r0 *1 0,2.775
X$1 3 5 1 2 6 SP6TCell
* cell instance $2 m0 *1 0,2.775
X$2 3 4 1 2 6 SP6TCell
.ENDS SP6TArray_2X1

* cell SP6TCell
* pin vdd
* pin wl
* pin bl
* pin bl_n
* pin vss
.SUBCKT SP6TCell 5 6 7 8 10
* net 5 vdd
* net 6 wl
* net 7 bl
* net 8 bl_n
* net 10 vss
* device instance $1 r0 *1 0.605,0.215 sky130_fd_pr__nfet_01v8__model
M$1 7 6 3 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.1113P
+ AD=0.18165P PS=1.37U PD=1.285U
* device instance $2 r0 *1 0.215,0.84 sky130_fd_pr__nfet_01v8__model
M$2 3 4 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.1113P PS=1.285U PD=1.37U
* device instance $3 r0 *1 1.575,0.215 sky130_fd_pr__nfet_01v8__model
M$3 8 6 4 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.1113P
+ AD=0.18165P PS=1.37U PD=1.285U
* device instance $4 r0 *1 1.965,0.84 sky130_fd_pr__nfet_01v8__model
M$4 4 3 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.42U AS=0.18165P
+ AD=0.1113P PS=1.285U PD=1.37U
* device instance $5 r0 *1 1.965,2.17 sky130_fd_pr__pfet_01v8__model
M$5 4 3 5 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1869P
+ AD=0.1113P PS=1.73U PD=1.37U
* device instance $6 r0 *1 0.215,2.17 sky130_fd_pr__pfet_01v8__model
M$6 5 4 3 5 sky130_fd_pr__pfet_01v8__model L=0.15U W=0.42U AS=0.1113P
+ AD=0.1869P PS=1.37U PD=1.73U
.ENDS SP6TCell
