.SUBCKT inv_chain 20 21
M$1 20 1 2 20 NCH_SVT_MAC L=0.016U W=3U 
M$2 20 2 3 20 NCH_SVT_MAC L=0.016U W=3U 
M$3 20 3 4 20 NCH_SVT_MAC L=0.016U W=3U 
M$4 20 4 5 20 NCH_SVT_MAC L=0.016U W=3U 
M$5 20 5 6 20 NCH_SVT_MAC L=0.016U W=3U 
M$6 20 6 7 20 NCH_SVT_MAC L=0.016U W=3U 
M$7 20 8 9 20 NCH_SVT_MAC L=0.016U W=3U 
M$8 20 9 10 20 NCH_SVT_MAC L=0.016U W=3U 
M$9 20 10 11 20 NCH_SVT_MAC L=0.016U W=3U 
M$10 20 11 12 20 NCH_SVT_MAC L=0.016U W=3U 
M$11 20 12 13 20 NCH_SVT_MAC L=0.016U W=3U 
M$12 20 14 15 20 NCH_SVT_MAC L=0.016U W=3U 
M$13 20 15 16 20 NCH_SVT_MAC L=0.016U W=3U 
M$14 20 16 17 20 NCH_SVT_MAC L=0.016U W=3U 
M$15 20 17 18 20 NCH_SVT_MAC L=0.016U W=3U 
M$16 20 18 19 20 NCH_SVT_MAC L=0.016U W=3U 
M$17 21 1 2 21 PCH_SVT_MAC L=0.016U W=3U 
M$18 21 2 3 21 PCH_SVT_MAC L=0.016U W=3U 
M$19 21 3 4 21 PCH_SVT_MAC L=0.016U W=3U 
M$20 21 4 5 21 PCH_SVT_MAC L=0.016U W=3U 
M$21 21 5 6 21 PCH_SVT_MAC L=0.016U W=3U 
M$22 21 6 7 21 PCH_SVT_MAC L=0.016U W=3U 
M$23 21 8 9 21 PCH_SVT_MAC L=0.016U W=3U 
M$24 21 9 10 21 PCH_SVT_MAC L=0.016U W=3U 
M$25 21 10 11 21 PCH_SVT_MAC L=0.016U W=3U 
M$26 21 11 12 21 PCH_SVT_MAC L=0.016U W=3U 
M$27 21 12 13 21 PCH_SVT_MAC L=0.016U W=3U 
M$28 21 14 15 21 PCH_SVT_MAC L=0.016U W=3U 
M$29 21 15 16 21 PCH_SVT_MAC L=0.016U W=3U 
M$30 21 16 17 21 PCH_SVT_MAC L=0.016U W=3U 
M$31 21 17 18 21 PCH_SVT_MAC L=0.016U W=3U 
M$32 21 18 19 21 PCH_SVT_MAC L=0.016U W=3U 
.ENDS inv_chain
