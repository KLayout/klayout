VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

LAYER M1
  TYPE ROUTING ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  WIDTH 0.05 ;
END M2

END LIBRARY
