magic
tech scmos
timestamp 1534324708
<< silk >>
rect 0 14 12 18
rect 8 11 12 14
rect 4 10 12 11
rect 1 8 12 10
rect 0 7 11 8
rect 0 4 4 7
rect 0 0 12 4
<< end >>
