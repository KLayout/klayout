VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

LAYER M1
  TYPE ROUTING ;
END M1
LAYER M2
  TYPE ROUTING ;
END M2

END LIBRARY
